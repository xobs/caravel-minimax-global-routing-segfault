* NGSPICE file created from minimax_rf.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

.subckt minimax_rf addrD[0] addrD[1] addrD[2] addrD[3] addrD[4] addrS[0] addrS[1]
+ addrS[2] addrS[3] addrS[4] clk new_value[0] new_value[10] new_value[11] new_value[12]
+ new_value[13] new_value[14] new_value[15] new_value[16] new_value[17] new_value[18]
+ new_value[19] new_value[1] new_value[20] new_value[21] new_value[22] new_value[23]
+ new_value[24] new_value[25] new_value[26] new_value[27] new_value[28] new_value[29]
+ new_value[2] new_value[30] new_value[31] new_value[3] new_value[4] new_value[5]
+ new_value[6] new_value[7] new_value[8] new_value[9] rD[0] rD[10] rD[11] rD[12] rD[13]
+ rD[14] rD[15] rD[16] rD[17] rD[18] rD[19] rD[1] rD[20] rD[21] rD[22] rD[23] rD[24]
+ rD[25] rD[26] rD[27] rD[28] rD[29] rD[2] rD[30] rD[31] rD[3] rD[4] rD[5] rD[6] rD[7]
+ rD[8] rD[9] rS[0] rS[10] rS[11] rS[12] rS[13] rS[14] rS[15] rS[16] rS[17] rS[18]
+ rS[19] rS[1] rS[20] rS[21] rS[22] rS[23] rS[24] rS[25] rS[26] rS[27] rS[28] rS[29]
+ rS[2] rS[30] rS[31] rS[3] rS[4] rS[5] rS[6] rS[7] rS[8] rS[9] vdd vss we
XANTENNA__12658__A2 register_file\[21\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09671_ _04913_ register_file\[27\]\[16\] _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11330__A2 _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08622_ _03808_ register_file\[26\]\[1\] _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09812__B _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08553_ _03879_ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15105__I _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11094__A1 _06064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08484_ _03810_ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07837__A2 register_file\[29\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12830__A2 _07377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09039__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14944__I _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14032__A1 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12594__A1 _07023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09105_ _04213_ register_file\[28\]\[7\] _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12464__I _07145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09036_ _04149_ register_file\[15\]\[6\] _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14335__A2 _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15532__A1 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12346__A1 _07016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12897__A2 register_file\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09938_ _05114_ register_file\[28\]\[20\] _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12649__A2 _07260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13846__A1 _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09514__A2 register_file\[8\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09869_ _05171_ _05177_ _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11900_ _06682_ _06792_ _06794_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12880_ _07406_ _07407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15891__CLK clknet_leaf_213_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11831_ _06748_ register_file\[7\]\[21\] _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12639__I _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13074__A2 _07520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15015__I _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14550_ _02058_ _02059_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11762_ _06708_ _06704_ _06709_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12821__A2 register_file\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13501_ _01021_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_41_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10713_ _03890_ register_file\[15\]\[31\] _06009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14481_ _01988_ _01991_ _01825_ _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__16247__CLK clknet_leaf_190_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14023__A1 _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11693_ _06650_ register_file\[8\]\[7\] _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16220_ _00608_ clknet_leaf_38_clk register_file\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13432_ _07737_ _07752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10644_ _05693_ register_file\[22\]\[30\] _05941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12585__A1 _07212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11388__A2 _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16151_ _00539_ clknet_leaf_190_clk register_file\[31\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13363_ _07553_ _07704_ _07710_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10575_ _05871_ _05872_ _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09450__A1 _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__A2 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15102_ _02604_ _02605_ _02276_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12314_ _07054_ register_file\[25\]\[9\] _07056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16397__CLK clknet_leaf_142_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10060__A2 register_file\[9\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14326__A2 register_file\[20\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15523__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16082_ _00470_ clknet_leaf_231_clk register_file\[4\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13294_ _07667_ register_file\[14\]\[24\] _07669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12337__A1 _07006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15033_ _02534_ _02536_ _02537_ _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12245_ _06112_ _07009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08005__A2 register_file\[31\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12176_ _06265_ _03815_ _06959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11560__A2 _06575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11127_ _06126_ _06300_ _06303_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11058_ _06218_ register_file\[28\]\[28\] _06261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15935_ _00323_ clknet_leaf_3_clk register_file\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10009_ _05114_ register_file\[20\]\[21\] _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15866_ _00254_ clknet_leaf_255_clk register_file\[12\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14817_ _02071_ register_file\[31\]\[14\] _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09269__A1 _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15797_ _00185_ clknet_leaf_205_clk register_file\[19\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11076__A1 _06033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14748_ _02169_ register_file\[20\]\[13\] _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12812__A2 _07360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10823__A1 _06100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14764__I _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14679_ _02103_ register_file\[10\]\[12\] _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16418_ _00806_ clknet_leaf_59_clk register_file\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_193_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15614__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12576__A1 _07212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12284__I _06163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16349_ _00737_ clknet_leaf_302_clk register_file\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10051__A2 register_file\[24\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09992__A2 register_file\[22\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15764__CLK clknet_leaf_177_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11000__A1 _06225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09744__A2 register_file\[24\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08547__A3 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07984_ _03235_ register_file\[21\]\[26\] _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13828__A1 _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09723_ _04830_ register_file\[10\]\[16\] _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11303__A2 _06408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09654_ _04962_ _04965_ _04900_ _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08937__I _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08605_ _03896_ _03931_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09585_ _04832_ register_file\[23\]\[14\] _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13056__A2 _07505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08158__B _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08536_ _03771_ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13999__B _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08467_ _03790_ _03792_ _03793_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__14005__A1 _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08398_ _03701_ register_file\[28\]\[31\] _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_5_31__f_clk_I clknet_3_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12567__A1 _06997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08235__A2 _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14308__A2 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15505__A1 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10360_ _05657_ _05660_ _04131_ _05661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12319__A1 _07054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09019_ _04054_ register_file\[11\]\[6\] _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11790__A2 _06720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10291_ _05527_ register_file\[23\]\[25\] _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12030_ _01532_ _06864_ _06872_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09735__A2 _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13819__A1 _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13981_ _01411_ register_file\[21\]\[4\] _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09499__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13295__A2 _07663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13753__I _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15720_ _00108_ clknet_leaf_88_clk register_file\[27\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12932_ _07417_ _07439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_98_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08847__I _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15651_ _00039_ clknet_leaf_53_clk register_file\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12369__I _07087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12863_ _07293_ _07391_ _07397_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14602_ _01693_ _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11058__A1 _06218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11814_ _06741_ register_file\[7\]\[14\] _06743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15582_ _03078_ _03079_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14795__A2 register_file\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15637__CLK clknet_leaf_211_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12794_ _07304_ _07350_ _07355_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14533_ _02043_ _01961_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11745_ _06696_ _06692_ _06697_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09671__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08474__A2 register_file\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14464_ _01972_ _01974_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11676_ _06647_ _06641_ _06648_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12558__A1 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16203_ _00591_ clknet_leaf_97_clk register_file\[24\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13415_ _07729_ _07742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10627_ _05922_ _05923_ _05924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14395_ _01650_ register_file\[31\]\[9\] _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16134_ _00522_ clknet_leaf_90_clk register_file\[31\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10033__A2 register_file\[29\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11230__A1 _06164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13346_ _07536_ _07697_ _07700_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09974__A2 register_file\[5\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10558_ _05731_ register_file\[8\]\[29\] _05856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11781__A2 _06720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16065_ _00453_ clknet_leaf_313_clk register_file\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13277_ _07653_ register_file\[14\]\[17\] _07659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10489_ _05589_ register_file\[20\]\[28\] _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_250_clk_I clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15016_ _02520_ register_file\[10\]\[16\] _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12228_ _06090_ _06997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12159_ _06701_ _06943_ _06949_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13286__A2 _07663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_265_clk_I clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15918_ _00306_ clknet_leaf_187_clk register_file\[10\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15027__A3 _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15849_ _00237_ clknet_leaf_111_clk register_file\[12\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13038__A2 _07458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10301__B _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11049__A1 _06254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09370_ _04413_ register_file\[9\]\[11\] _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14786__A2 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12797__A1 _07311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08321_ _03352_ register_file\[10\]\[30\] _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08252_ _01048_ register_file\[13\]\[29\] _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10272__A2 _05573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_203_clk_I clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12549__A1 _07190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ _03512_ _03361_ _03513_ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_158_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13210__A2 _07615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10024__A2 register_file\[4\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11221__A1 _06355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_218_clk_I clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14710__A2 register_file\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11524__A2 _06554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10262__I _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12898__B _07419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input36_I new_value[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07967_ _03300_ _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14474__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13573__I _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16092__CLK clknet_leaf_301_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09706_ _04750_ register_file\[19\]\[16\] _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07898_ _03228_ _03230_ _03231_ _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ _04750_ register_file\[7\]\[15\] _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12189__I _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14226__A1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10211__B _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07900__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09568_ _04750_ register_file\[11\]\[14\] _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12788__A1 _07298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08519_ _03842_ _03845_ _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09499_ _04812_ register_file\[4\]\[13\] _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09498__I _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11460__A1 _06517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11530_ _06558_ register_file\[11\]\[9\] _06560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10263__A2 register_file\[28\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09405__A1 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11461_ _06402_ _06513_ _06518_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13201__A2 _07608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13200_ _07612_ register_file\[15\]\[18\] _07613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10015__A2 register_file\[17\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11212__A1 _06355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10412_ _05699_ _05712_ _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11392_ _06476_ register_file\[26\]\[18\] _06477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09956__A2 register_file\[8\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14180_ _01605_ register_file\[15\]\[6\] _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13748__I register_file\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13131_ _07563_ register_file\[16\]\[25\] _07569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09447__B _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10343_ _05636_ _05644_ _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13062_ _07519_ _07520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10274_ _05571_ _05576_ _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12712__A1 _07304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16435__CLK clknet_leaf_167_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12013_ _06815_ register_file\[5\]\[31\] _06861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09961__I _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13483__I _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11279__A1 _06400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10900__I _06163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13964_ _01216_ register_file\[31\]\[4\] _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16585__CLK clknet_leaf_114_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__A1 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15703_ _00091_ clknet_leaf_212_clk register_file\[28\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12915_ _07409_ _07429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12099__I _06913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09892__A1 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13895_ _01409_ _01410_ _01412_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_61_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15634_ _00022_ clknet_leaf_178_clk register_file\[30\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12846_ _07276_ _07384_ _07387_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15565_ _01068_ _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12777_ _07340_ register_file\[20\]\[22\] _07346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09644__A1 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08447__A2 register_file\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15203__I register_file\[4\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14516_ _01142_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11451__A1 _06393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11728_ _06684_ _06680_ _06685_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15496_ _02992_ _02994_ _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14447_ _01956_ _01958_ _01709_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15193__A2 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11659_ _06591_ register_file\[10\]\[30\] _06636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11203__A1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14940__A2 _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14378_ _01849_ _01890_ _01634_ net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13658__I _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16117_ _00505_ clknet_leaf_221_clk register_file\[3\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12951__A1 _07407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13329_ _07686_ register_file\[29\]\[5\] _07691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_1_0_clk clknet_0_clk clknet_3_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16048_ _00436_ clknet_leaf_230_clk register_file\[5\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12703__A1 _07298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ _04184_ _04192_ _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07821_ _02903_ register_file\[23\]\[24\] _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13259__A2 _07642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10190__A1 _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13393__I _07727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_84_clk_I clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10810__I _06090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09092__B _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08487__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08135__A1 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14208__A1 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09883__A1 _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10031__B _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15952__CLK clknet_leaf_216_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09422_ _04669_ register_file\[20\]\[12\] _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11690__A1 _06650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14759__A2 register_file\[8\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_99_clk_I clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09353_ _03843_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13431__A2 _07745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_142_clk_I clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08304_ _03631_ _03632_ _01126_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11442__A1 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09284_ _04600_ register_file\[18\]\[10\] _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_clk_I clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11993__A2 register_file\[5\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08235_ _03563_ _01133_ _03564_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13195__A1 _07605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09938__A2 register_file\[28\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08166_ _03493_ _03496_ _03340_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_157_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07949__A1 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12942__A1 _07443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11745__A2 _06692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16458__CLK clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08097_ _03428_ _03102_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_37_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08374__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15239__A3 _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12170__A2 _06950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08999_ _04319_ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11816__I _06729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14998__A2 register_file\[21\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08126__A1 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10961_ _06196_ register_file\[2\]\[22\] _06202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12700_ _07295_ _07296_ _07297_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13680_ _01200_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_71_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10892_ _06156_ _06140_ _06157_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12631_ _07242_ register_file\[21\]\[5\] _07249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12647__I _07247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09626__A1 _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13422__A2 _07745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11551__I _06542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15350_ _02520_ register_file\[10\]\[20\] _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10236__A2 register_file\[13\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11433__A1 _06375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12562_ _06992_ _07201_ _07204_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_169_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14301_ _01813_ register_file\[27\]\[8\] _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11984__A2 register_file\[5\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11513_ _06375_ _06544_ _06549_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15281_ register_file\[7\]\[19\] _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12493_ _07157_ register_file\[23\]\[17\] _07163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15175__A2 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13186__A1 _07536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14232_ _01068_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09929__A2 register_file\[2\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11444_ _06386_ _06506_ _06508_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08860__I _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12933__A1 _07436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13478__I _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14163_ _01675_ _01677_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11375_ _06462_ register_file\[26\]\[11\] _06467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13114_ _07551_ register_file\[16\]\[20\] _07557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10326_ _05624_ _05627_ _03795_ _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14094_ _01599_ _01609_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13045_ _07507_ register_file\[16\]\[0\] _07508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10257_ _05558_ _05559_ _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09691__I _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08365__A1 _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10188_ _05490_ _05491_ _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10172__A1 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14438__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11726__I _06103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15975__CLK clknet_leaf_297_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14102__I register_file\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14996_ _02497_ _02500_ _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14989__A2 register_file\[17\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08117__A1 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13110__A1 _07551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13947_ _01202_ register_file\[24\]\[4\] _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09865__A1 _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08668__A2 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11672__A1 _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10475__A2 register_file\[1\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13878_ _01390_ _01393_ _01395_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15617_ _00005_ clknet_leaf_19_clk register_file\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12829_ _07374_ register_file\[1\]\[10\] _07378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16597_ _00985_ clknet_leaf_217_clk register_file\[9\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15548_ _02964_ register_file\[2\]\[22\] _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_187_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11975__A2 _06833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_150_clk clknet_5_30__leaf_clk clknet_leaf_150_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15479_ _01009_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08840__A2 register_file\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16600__CLK clknet_leaf_257_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13177__A1 _07526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08020_ _03352_ register_file\[10\]\[26\] _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08770__I _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12924__A1 _07274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11727__A2 register_file\[8\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10805__I _06028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09971_ _05272_ _05277_ _04191_ _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08922_ _04242_ _04243_ _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12152__A2 _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08853_ _04166_ _04175_ _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11636__I _06601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07804_ _03098_ _03139_ _02888_ net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08784_ _03956_ register_file\[22\]\[3\] _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08108__A1 _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13101__A1 _07546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13851__I _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10466__A2 register_file\[25\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16130__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09405_ _04582_ register_file\[28\]\[12\] _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09608__A1 _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14601__A1 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13404__A2 _07728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09336_ _04516_ register_file\[6\]\[11\] _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11415__A1 _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11966__A2 _06833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09267_ _04581_ _04583_ _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16280__CLK clknet_leaf_191_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_141_clk clknet_5_26__leaf_clk clknet_leaf_141_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_107_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08831__A2 register_file\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08218_ _03546_ _01084_ _03547_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09198_ _03807_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11718__A2 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08149_ _03476_ _03479_ _01101_ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11160_ _06322_ register_file\[13\]\[2\] _06325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14668__A1 _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14631__B _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10111_ _03847_ _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11091_ _06060_ _06279_ _06282_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08347__A1 _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10042_ _05328_ _05347_ _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output67_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10154__A1 _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13891__A2 register_file\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10450__I _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14850_ _02355_ _02356_ _02276_ _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13801_ _01319_ register_file\[28\]\[2\] _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14781_ _02288_ _02203_ _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09847__A1 _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11993_ _06844_ register_file\[5\]\[22\] _06850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16520_ _00908_ clknet_leaf_46_clk register_file\[14\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13732_ _01246_ _01251_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10944_ _06177_ _06192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10457__A2 register_file\[29\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11654__A1 _06436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16451_ _00839_ clknet_leaf_56_clk register_file\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13663_ _01177_ _01180_ _01183_ _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15396__A2 register_file\[18\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11281__I _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10875_ _06143_ _06144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15402_ _02736_ register_file\[22\]\[21\] _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11406__A1 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12614_ _07230_ _07233_ _07236_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16382_ _00770_ clknet_leaf_29_clk register_file\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09075__A2 register_file\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13594_ _01114_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15333_ _02832_ _02833_ _02751_ _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11957__A2 register_file\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12545_ _07190_ register_file\[22\]\[5\] _07195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_132_clk clknet_5_26__leaf_clk clknet_leaf_132_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13159__A1 _07509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15264_ _02513_ register_file\[9\]\[19\] _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08590__I _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12476_ _07145_ _07153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_145_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12906__A1 _07422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14215_ _01557_ register_file\[26\]\[7\] _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11427_ _06497_ _06498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15195_ _02444_ register_file\[15\]\[18\] _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12382__A2 _07088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14146_ _01405_ register_file\[18\]\[6\] _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11358_ _06380_ _06448_ _06456_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10393__A1 _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16003__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13936__I register_file\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12840__I _07369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10309_ _05608_ _05610_ _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15320__A2 register_file\[30\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14077_ _01591_ _01592_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11289_ _06403_ register_file\[19\]\[15\] _06409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08338__A1 _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13331__A1 _07686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13028_ _07298_ _07494_ _07496_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_199_clk clknet_5_19__leaf_clk clknet_leaf_199_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08889__A2 register_file\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11893__A1 _06674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15084__A1 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16153__CLK clknet_leaf_191_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09838__A1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14979_ _02235_ register_file\[28\]\[16\] _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11645__A1 _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13398__A1 _07730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09066__A2 register_file\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09121_ _04438_ _04439_ _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11948__A2 _06816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15139__A2 register_file\[17\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_123_clk clknet_5_24__leaf_clk clknet_leaf_123_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_175_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08813__A2 register_file\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09052_ _04090_ register_file\[14\]\[7\] _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14898__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08003_ _03334_ _03089_ _03335_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12373__A2 _07088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13570__A1 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09954_ _05251_ _05260_ _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09545__B _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08329__A1 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07844__I _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08905_ _04210_ _04227_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09885_ _05192_ register_file\[27\]\[19\] _05193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10136__A1 _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ _04141_ _04159_ _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08767_ _04090_ register_file\[14\]\[3\] _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09829__A1 _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14822__A1 _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10439__A2 register_file\[12\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08675__I _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08698_ _03808_ register_file\[22\]\[2\] _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12197__I _06962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output105_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13389__A1 _07679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10660_ _05956_ _03928_ _05957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09057__A2 register_file\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14050__A2 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14626__B _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09319_ _03927_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_107_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12061__A1 _06885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_114_clk clknet_5_13__leaf_clk clknet_leaf_114_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10591_ _03887_ register_file\[6\]\[29\] _05889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08804__A2 register_file\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12330_ _06999_ _07064_ _07065_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_194_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10611__A2 register_file\[24\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16026__CLK clknet_leaf_252_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12261_ _07018_ _07012_ _07020_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15550__A2 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14000_ _01513_ _01516_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11212_ _06355_ register_file\[13\]\[23\] _06356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12364__A2 _07042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13561__A1 _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12192_ _06969_ _06961_ _06971_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12660__I _06090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput53 net53 rD[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11143_ _06156_ _06307_ _06312_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09455__B _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput64 net64 rD[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput75 net75 rD[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_150_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput86 net86 rS[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__12116__A2 _06922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput97 net97 rS[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_150_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15951_ _00339_ clknet_leaf_189_clk register_file\[8\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10127__A1 _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11074_ _06021_ _06269_ _06272_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14902_ _02406_ _02323_ _02407_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10025_ _05329_ _05330_ _05331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15882_ _00270_ clknet_leaf_112_clk register_file\[11\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10678__A2 register_file\[29\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15066__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08740__A1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14833_ _02258_ register_file\[21\]\[14\] _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13616__A2 _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11627__A1 _06613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14764_ _01426_ _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11976_ _06825_ _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_63_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13715_ _01097_ register_file\[31\]\[1\] _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16503_ _00891_ clknet_leaf_222_clk register_file\[15\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10927_ _06169_ _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14695_ _02202_ _02203_ _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16434_ _00822_ clknet_leaf_165_clk register_file\[17\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13646_ _01166_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10850__A2 _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09048__A2 register_file\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10858_ _06129_ _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12835__I _07361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16365_ _00753_ clknet_leaf_143_clk register_file\[1\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12052__A1 _06885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_105_clk clknet_5_15__leaf_clk clknet_leaf_105_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13577_ _01097_ register_file\[31\]\[0\] _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10789_ _06051_ _06074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_125_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15316_ _02651_ register_file\[28\]\[20\] _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12528_ _07182_ _07183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_5_17__f_clk clknet_3_4_0_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16296_ _00684_ clknet_leaf_80_clk register_file\[21\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15247_ _02581_ register_file\[27\]\[19\] _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12459_ _07142_ register_file\[23\]\[3\] _07143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12355__A2 register_file\[25\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13552__A1 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16519__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15178_ _02660_ _02680_ _02347_ _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_5_8__f_clk_I clknet_3_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09220__A2 _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10366__A1 _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13666__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14129_ _01640_ _01643_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12107__A2 register_file\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13304__A1 _07574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07782__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10090__I _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09670_ _04781_ register_file\[26\]\[16\] _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08621_ _03945_ _03946_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11618__A1 _06400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08552_ _03764_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15693__CLK clknet_leaf_148_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11094__A2 _06279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08483_ _03784_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_74_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16049__CLK clknet_leaf_230_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09104_ _04211_ register_file\[29\]\[7\] _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12594__A2 _07222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08262__A3 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09035_ _04146_ register_file\[14\]\[6\] _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15532__A2 register_file\[15\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16199__CLK clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12346__A2 _07071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10357__A1 _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13576__I _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15296__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08970__A1 _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09937_ _05112_ register_file\[29\]\[20\] _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10109__A1 _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09868_ _05176_ _04973_ _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15048__A1 _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08819_ _03901_ register_file\[4\]\[3\] _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15599__A2 _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09799_ _05108_ _04973_ _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11609__A1 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14200__I register_file\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11830_ _06691_ _06751_ _06752_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12282__A1 _06960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11761_ _06699_ register_file\[8\]\[27\] _06709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13500_ net8 _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_41_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10712_ _03887_ register_file\[14\]\[31\] _06008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14480_ _01989_ _01906_ _01990_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11692_ _06059_ _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15220__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14023__A2 register_file\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13431_ _07541_ _07745_ _07751_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10643_ _05938_ _05939_ _05940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__A1 _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12585__A2 register_file\[22\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16150_ _00538_ clknet_leaf_181_clk register_file\[31\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13782__A1 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13362_ _07708_ register_file\[29\]\[19\] _07710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10574_ _03844_ register_file\[24\]\[29\] _05872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10596__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15101_ _02520_ register_file\[10\]\[17\] _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12313_ _06982_ _07050_ _07055_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16081_ _00469_ clknet_5_21__leaf_clk register_file\[4\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13293_ _07562_ _07663_ _07668_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12337__A2 _07064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15032_ _01158_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12244_ _07006_ _07000_ _07008_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10348__A1 _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12175_ _06020_ _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11126_ _06297_ register_file\[27\]\[22\] _06303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13837__A2 _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11057_ _06148_ _06257_ _06260_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11848__A1 _06710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15934_ _00322_ clknet_leaf_305_clk register_file\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10008_ _05112_ register_file\[21\]\[21\] _05314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10520__A1 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15865_ _00253_ clknet_leaf_260_clk register_file\[12\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14816_ _01045_ _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09269__A2 register_file\[23\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15796_ _00184_ clknet_leaf_172_clk register_file\[19\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12273__A1 _07019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11076__A2 _06269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14747_ _02250_ _02254_ _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11959_ _06817_ _06830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10823__A2 _06096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14678_ _02101_ register_file\[11\]\[12\] _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16417_ _00805_ clknet_leaf_59_clk register_file\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13629_ _01128_ _01149_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12576__A2 register_file\[22\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16348_ _00736_ clknet_leaf_281_clk register_file\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16279_ _00667_ clknet_leaf_197_clk register_file\[22\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15514__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10339__A1 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16491__CLK clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10813__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11000__A2 register_file\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08952__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07983_ _03068_ register_file\[20\]\[26\] _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13828__A2 register_file\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09722_ _05031_ _05032_ _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11839__A1 _06701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09653_ _04963_ _04964_ _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10511__A1 _05794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15116__I _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08604_ _03915_ _03930_ _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08180__A2 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09584_ _04830_ register_file\[22\]\[14\] _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15450__A1 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14253__A2 _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08535_ _03861_ register_file\[13\]\[0\] _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12264__A1 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08466_ net3 _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_195_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08397_ _03722_ _03724_ _01094_ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12567__A2 _07201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15505__A2 register_file\[28\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12319__A2 register_file\[25\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09018_ _04052_ register_file\[10\]\[6\] _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10290_ _05525_ register_file\[22\]\[25\] _05592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09196__A1 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15269__A1 _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13980_ _01319_ register_file\[20\]\[4\] _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12931_ _07281_ _07432_ _07438_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16214__CLK clknet_leaf_207_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15650_ _00038_ clknet_5_8__leaf_clk register_file\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12862_ _07395_ register_file\[1\]\[24\] _07397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15441__A1 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14601_ _02025_ register_file\[14\]\[11\] _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11813_ _06674_ _06737_ _06742_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15581_ _02993_ register_file\[17\]\[23\] _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12793_ _07311_ register_file\[20\]\[29\] _07355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09120__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14532_ _02037_ _02042_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11744_ _06687_ register_file\[8\]\[22\] _06697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16364__CLK clknet_leaf_140_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09671__A2 register_file\[27\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14463_ _01973_ register_file\[25\]\[10\] _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12007__A1 _06815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11675_ _06643_ register_file\[8\]\[2\] _06648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12558__A2 _07201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16202_ _00590_ clknet_leaf_96_clk register_file\[24\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13414_ _07524_ _07738_ _07741_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10626_ _05674_ register_file\[16\]\[30\] _05923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14394_ _01045_ _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16133_ _00521_ clknet_leaf_79_clk register_file\[31\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13345_ _07694_ register_file\[29\]\[12\] _07700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11230__A2 _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ _05729_ register_file\[9\]\[29\] _05855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07985__A2 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16064_ _00452_ clknet_5_1__leaf_clk register_file\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13276_ _07546_ _07656_ _07658_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10488_ _05587_ register_file\[21\]\[28\] _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09187__A1 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15015_ _01138_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11729__I _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12227_ _06994_ _06988_ _06996_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14180__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12158_ _06947_ register_file\[3\]\[24\] _06949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10741__A1 _06033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11109_ _06278_ _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_116_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12089_ _06863_ net32 _06907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07942__I _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15917_ _00305_ clknet_leaf_121_clk register_file\[10\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12494__A1 _07004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11464__I _06505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08162__A2 _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15848_ _00236_ clknet_leaf_108_clk register_file\[12\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12246__A1 _07007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11049__A2 register_file\[28\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15779_ _00167_ clknet_leaf_56_clk register_file\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09111__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08320_ _03350_ register_file\[11\]\[30\] _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09662__A2 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08251_ _03356_ register_file\[12\]\[29\] _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10808__I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15731__CLK clknet_leaf_177_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08182_ _03276_ register_file\[15\]\[28\] _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11221__A2 register_file\[13\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15881__CLK clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10980__A1 _06160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08925__A1 _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16237__CLK clknet_leaf_139_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09553__B _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07966_ _03298_ _03299_ _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14474__A2 register_file\[28\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09705_ _04748_ register_file\[18\]\[16\] _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input29_I new_value[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12485__A1 _06994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07897_ _01559_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_94_clk clknet_5_14__leaf_clk clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09350__A1 _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09636_ _04748_ register_file\[6\]\[15\] _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16387__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14226__A2 register_file\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07900__A2 register_file\[28\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12237__A1 _07002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09567_ _04748_ register_file\[10\]\[14\] _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14777__A3 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12788__A2 _07350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08518_ _03844_ register_file\[16\]\[0\] _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09498_ _04124_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_23_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_310_clk_I clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08449_ _03762_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13737__A1 _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11460_ _06517_ register_file\[12\]\[13\] _06518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09405__A2 register_file\[28\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10411_ _05706_ _05711_ _05712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11212__A2 register_file\[13\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11391_ _06446_ _06476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output97_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13130_ _07519_ _07568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10342_ _05642_ _05643_ _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10971__A1 _06203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14162__A1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13061_ _07506_ _07519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10273_ _05575_ _05309_ _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14701__A3 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08916__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12012_ _06714_ _06818_ _06860_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12712__A2 _07296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10723__A1 _05989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09463__B _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11279__A2 _06396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13963_ _01045_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11284__I _06090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_85_clk clknet_5_11__leaf_clk clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08144__A2 register_file\[29\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15702_ _00090_ clknet_leaf_212_clk register_file\[28\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12914_ _07264_ _07425_ _07428_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13894_ _01411_ register_file\[29\]\[3\] _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15414__A1 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12845_ _07381_ register_file\[1\]\[17\] _07387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15633_ _00021_ clknet_leaf_165_clk register_file\[30\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08593__I _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13976__A1 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12776_ _07286_ _07343_ _07345_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15564_ _03061_ _01066_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09644__A2 register_file\[31\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14515_ _02025_ register_file\[14\]\[10\] _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11727_ _06675_ register_file\[8\]\[17\] _06685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15495_ _02993_ register_file\[25\]\[22\] _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11451__A2 _06506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13728__A1 _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14446_ _01957_ _01707_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11658_ _06440_ _06630_ _06635_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10609_ _05902_ _05905_ _04037_ _05906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12400__A1 _06990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11203__A2 _06344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14377_ _01869_ _01889_ _01632_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11589_ _06366_ _06592_ _06595_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16116_ _00504_ clknet_leaf_221_clk register_file\[3\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13328_ _07689_ _07690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08080__A1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10962__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11459__I _06497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14153__A1 _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13259_ _07529_ _07642_ _07648_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16047_ _00435_ clknet_leaf_245_clk register_file\[5\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08907__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12703__A2 _07296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13674__I _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09580__A1 _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07820_ _01325_ _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10190__A2 register_file\[15\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12467__A1 _07142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_76_clk clknet_5_10__leaf_clk clknet_leaf_76_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08135__A2 register_file\[25\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09421_ _04667_ register_file\[21\]\[12\] _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12219__A1 _06983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07894__A1 _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11690__A2 register_file\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09352_ _04667_ register_file\[29\]\[11\] _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13967__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08303_ _01090_ register_file\[26\]\[30\] _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09283_ _03904_ _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11442__A2 _06506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08234_ _01135_ register_file\[29\]\[29\] _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08165_ _03494_ _01141_ _03495_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_146_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12942__A2 register_file\[18\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08071__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08096_ _03426_ _03427_ _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10953__A1 _06108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15627__CLK clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14695__A2 _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10705__A1 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13584__I _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__A1 _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08374__A2 register_file\[8\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08998_ _03830_ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_75_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07949_ _03282_ register_file\[6\]\[25\] _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_47_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_67_clk clknet_5_10__leaf_clk clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__15777__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10960_ _06122_ _06199_ _06201_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11130__A1 _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09619_ _04663_ register_file\[15\]\[15\] _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07885__A1 _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10891_ _06026_ register_file\[30\]\[29\] _06157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15304__I _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12630_ _07247_ _07248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09626__A2 register_file\[10\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08429__A3 _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12561_ _07198_ register_file\[22\]\[12\] _07204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11433__A2 _06496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14300_ _01014_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11512_ _06546_ register_file\[11\]\[2\] _06549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15280_ _02450_ register_file\[6\]\[19\] _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_19_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12492_ _07002_ _07160_ _07162_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14231_ _01744_ _01490_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_264_clk_I clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12663__I _06094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13186__A2 _07601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11443_ _06502_ register_file\[12\]\[6\] _06508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16402__CLK clknet_leaf_159_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11197__A1 _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12933__A2 register_file\[18\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14162_ _01676_ register_file\[9\]\[6\] _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11374_ _06395_ _06465_ _06466_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13113_ _07519_ _07556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10325_ _05625_ _05626_ _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14093_ _01602_ _01607_ _01608_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14686__A2 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_279_clk_I clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13044_ _07506_ _07507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16552__CLK clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10256_ _05361_ register_file\[27\]\[24\] _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13494__I _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09562__A1 _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08365__A2 register_file\[3\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10187_ _05425_ register_file\[12\]\[23\] _05491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10172__A2 register_file\[27\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_202_clk_I clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14995_ _02498_ _02499_ _02336_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_58_clk clknet_5_8__leaf_clk clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09314__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13946_ _01419_ _01463_ _01201_ net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14539__B _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13877_ _01394_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11672__A2 register_file\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_217_clk_I clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15616_ _00004_ clknet_leaf_19_clk register_file\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12828_ _07369_ _07377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_22_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16596_ _00984_ clknet_leaf_214_clk register_file\[9\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15547_ _03045_ _02793_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12759_ _07269_ _07329_ _07335_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15478_ _02976_ _02808_ _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13177__A2 _07594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16082__CLK clknet_leaf_231_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14429_ _01937_ _01940_ _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11188__A1 _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12924__A2 _07432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10935__A1 _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14126__A1 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09970_ _05274_ _05276_ _05277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09882__I _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14677__A2 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08921_ _04172_ register_file\[19\]\[5\] _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12688__A1 _07279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08356__A2 _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10821__I _06099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08852_ _04169_ _04174_ _04102_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07803_ _03118_ _03138_ _02886_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08783_ _04105_ _04106_ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_49_clk clknet_5_9__leaf_clk clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08108__A2 register_file\[15\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09305__A1 _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13101__A2 _07544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11112__A1 _06290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12748__I _07321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12860__A1 _07395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09404_ _04580_ register_file\[29\]\[12\] _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09122__I _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14601__A2 register_file\[14\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09335_ _04649_ _04650_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11415__A2 register_file\[26\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16425__CLK clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09266_ _04582_ register_file\[20\]\[10\] _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08292__A1 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13579__I _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08217_ _03235_ register_file\[21\]\[29\] _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12483__I _07137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09197_ _04513_ _04514_ _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11179__A1 _06069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08148_ _03477_ _03155_ _03478_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16575__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10926__A1 _06060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09792__A1 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ _03410_ _02912_ _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14668__A2 register_file\[23\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10110_ _05413_ _05414_ _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12679__A1 _07281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11090_ _06275_ register_file\[27\]\[7\] _06282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10041_ _05337_ _05346_ _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10731__I _06025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10154__A2 register_file\[16\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11351__A1 _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13800_ _01318_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11103__A1 _06082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14780_ register_file\[7\]\[13\] _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11992_ _06694_ _06847_ _06849_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10943_ _06091_ _06185_ _06191_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13731_ _01248_ _01250_ _01126_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12851__A1 _07281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11654__A2 _06630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16450_ _00838_ clknet_leaf_52_clk register_file\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10874_ _06142_ _06143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13662_ _01181_ _01182_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_3_0_0_clk clknet_0_clk clknet_3_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_108_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15401_ _02899_ _02733_ _02900_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12613_ _07235_ register_file\[21\]\[0\] _07236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11406__A2 register_file\[26\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12603__A1 _07183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16381_ _00769_ clknet_leaf_29_clk register_file\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13593_ _01004_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12544_ _07193_ _07194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15332_ _02667_ register_file\[18\]\[20\] _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08283__A1 _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13489__I _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14356__A1 _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13159__A2 _07584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12475_ _06985_ _07146_ _07152_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_83_clk_I clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15263_ _02764_ register_file\[8\]\[19\] _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10906__I _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12906__A2 register_file\[18\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11426_ _06494_ _06497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14214_ _01382_ register_file\[27\]\[7\] _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15194_ _02442_ register_file\[14\]\[18\] _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10917__A1 _06174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14108__A1 _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09783__A1 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14145_ _01313_ register_file\[19\]\[6\] _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11357_ _06454_ register_file\[26\]\[4\] _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15942__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11590__A1 _06594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10308_ _05609_ register_file\[15\]\[25\] _05610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_98_clk_I clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14076_ _01242_ register_file\[9\]\[5\] _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11288_ _06383_ _06408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11737__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13027_ _07491_ register_file\[17\]\[26\] _07496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_141_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _05273_ register_file\[14\]\[24\] _05542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13331__A2 register_file\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11342__A1 _06444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15608__A1 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11893__A2 _06785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15084__A2 register_file\[21\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14978_ _02479_ _02482_ _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_156_clk_I clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12568__I _07193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12842__A1 _07271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13929_ _01162_ _01446_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11645__A2 _06623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16448__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_36_clk_I clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13398__A2 register_file\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16579_ _00967_ clknet_leaf_13_clk register_file\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09120_ _04369_ register_file\[28\]\[8\] _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08274__A1 _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12070__A2 _06895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16598__CLK clknet_leaf_224_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10081__A1 _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09051_ _04368_ _04370_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10816__I _06051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08002_ _03090_ register_file\[29\]\[26\] _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10908__A1 _06170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11581__A1 _06543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09953_ _05256_ _05259_ _04452_ _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_109_clk_I clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08904_ _04221_ _04226_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09884_ _03810_ _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10136__A2 register_file\[3\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11333__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08835_ _04152_ _04158_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15075__A2 _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13086__A1 _07527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09561__B _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08766_ _03779_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09829__A2 register_file\[8\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input11_I new_value[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14822__A2 register_file\[17\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_25__f_clk_I clknet_3_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12833__A1 _07374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08697_ _04020_ _04021_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15815__CLK clknet_leaf_107_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14693__I register_file\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13389__A2 register_file\[29\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09318_ _04631_ _04632_ _04634_ _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12061__A2 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10590_ _05886_ _05887_ _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14338__A1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09249_ _04291_ register_file\[1\]\[9\] _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10726__I _06020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15965__CLK clknet_leaf_307_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14889__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12260_ _07019_ register_file\[31\]\[23\] _07020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13010__A1 _07484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11211_ _06318_ _06355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12191_ _06970_ register_file\[31\]\[3\] _06971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11572__A1 _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11142_ _06268_ register_file\[27\]\[29\] _06312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput54 net54 rD[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_150_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput65 net65 rD[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_122_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09517__A1 _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput76 net76 rS[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput87 net87 rS[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_153_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15950_ _00338_ clknet_leaf_189_clk register_file\[8\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11073_ _06271_ register_file\[27\]\[0\] _06272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput98 net98 rS[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_62_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11324__A1 _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09027__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14901_ _02071_ register_file\[31\]\[15\] _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10024_ _05063_ register_file\[4\]\[21\] _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15881_ _00269_ clknet_5_13__leaf_clk register_file\[11\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11875__A2 register_file\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15066__A2 register_file\[30\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14832_ _02169_ register_file\[20\]\[14\] _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09471__B _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13077__A1 _07529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14813__A2 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12824__A1 _07374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14763_ _02269_ _02270_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11975_ _06677_ _06833_ _06839_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16502_ _00890_ clknet_leaf_225_clk register_file\[15\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13714_ _01090_ register_file\[30\]\[1\] _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10926_ _06060_ _06178_ _06181_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14694_ _01354_ _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16433_ _00821_ clknet_leaf_162_clk register_file\[17\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13645_ _00998_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10857_ _06128_ _06129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16364_ _00752_ clknet_leaf_140_clk register_file\[1\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10788_ _06072_ _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13576_ _01096_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12052__A2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10063__A1 _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14329__A1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15315_ _02810_ _02815_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12527_ _06023_ _03991_ _07182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16295_ _00683_ clknet_leaf_80_clk register_file\[21\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13012__I _07465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13001__A1 _07477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15246_ _02747_ _01225_ _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12458_ _07137_ _07142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09756__A1 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11409_ _06483_ register_file\[26\]\[25\] _06487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13552__A2 register_file\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12389_ _07094_ register_file\[24\]\[7\] _07101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09646__B _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15177_ _02670_ _02679_ _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10366__A2 register_file\[6\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07945__I _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16120__CLK clknet_leaf_241_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14128_ _01641_ _01642_ _01560_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09508__A1 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10371__I _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13304__A2 _07670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14059_ _01573_ _01574_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input3_I addrD[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16270__CLK clknet_leaf_153_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15057__A2 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13682__I _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08620_ _03803_ register_file\[24\]\[1\] _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14804__A2 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08551_ _03866_ _03873_ _03877_ _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12298__I _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11618__A2 _06609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08482_ _03808_ register_file\[30\]\[0\] _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08495__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15988__CLK clknet_leaf_229_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08247__A1 _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12043__A2 _06874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13240__A1 _07634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09103_ _04412_ _04422_ _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10054__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09034_ _04353_ _04354_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09747__A1 _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13543__A2 _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11554__A1 _06572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10357__A2 register_file\[26\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14099__A3 _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08970__A2 register_file\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_280_clk clknet_5_6__leaf_clk clknet_leaf_280_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10281__I _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09936_ _05212_ _05243_ _04977_ net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_154_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11306__A1 _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09867_ _05172_ _05174_ _05175_ _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15048__A2 register_file\[1\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08818_ _03898_ register_file\[5\]\[3\] _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13059__A1 _07516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07804__B _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09798_ _05105_ _05106_ _05107_ _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11609__A2 _06602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08749_ _03905_ register_file\[30\]\[2\] _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12806__A1 _07362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_23__f_clk clknet_3_5_0_clk clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11760_ _06147_ _06708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12282__A2 register_file\[31\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10711_ _06005_ _06006_ _06007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11691_ _06658_ _06656_ _06659_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11840__I _06729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13430_ _07749_ register_file\[9\]\[14\] _07751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10642_ _05758_ register_file\[20\]\[30\] _05939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12034__A2 _06874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13361_ _07550_ _07704_ _07709_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10456__I _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08789__A2 register_file\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10573_ _03841_ register_file\[25\]\[29\] _05871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13782__A2 register_file\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15100_ _02518_ register_file\[11\]\[17\] _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11793__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10596__A2 register_file\[3\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12312_ _07054_ register_file\[25\]\[8\] _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16143__CLK clknet_leaf_153_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13292_ _07667_ register_file\[14\]\[23\] _07668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16080_ _00468_ clknet_leaf_234_clk register_file\[4\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12243_ _07007_ register_file\[31\]\[18\] _07008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15031_ _02535_ _02203_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14731__A1 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11545__A1 _06565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10348__A2 register_file\[16\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12174_ _06716_ _06914_ _06957_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11287__I _06094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10405__B _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16293__CLK clknet_leaf_75_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11125_ _06122_ _06300_ _06302_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_271_clk clknet_5_7__leaf_clk clknet_leaf_271_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13298__A1 _07567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11056_ _06254_ register_file\[28\]\[27\] _06260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15933_ _00321_ clknet_leaf_307_clk register_file\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11848__A2 _06758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10007_ _05280_ _05312_ _05313_ net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08596__I _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15864_ _00252_ clknet_leaf_260_clk register_file\[12\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14815_ _02321_ register_file\[30\]\[14\] _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14798__A1 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15795_ _00183_ clknet_leaf_172_clk register_file\[19\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13007__I _07454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14746_ _02251_ _02253_ _01919_ _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08477__A1 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12273__A2 register_file\[31\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11958_ _06660_ _06826_ _06829_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13470__A1 _07580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10909_ _06021_ _06168_ _06171_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14677_ _02185_ _01855_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11889_ _06782_ register_file\[6\]\[12\] _06788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11750__I _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16416_ _00804_ clknet_leaf_15_clk register_file\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08229__A1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13628_ _01137_ _01145_ _01148_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12025__A2 _06864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13222__A1 _07572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09977__A1 _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14970__A1 _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16347_ _00735_ clknet_leaf_272_clk register_file\[20\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13559_ _01079_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11784__A1 _06722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10587__A2 _05884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16278_ _00666_ clknet_leaf_207_clk register_file\[22\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15514__A3 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13677__I _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09729__A1 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15229_ _02727_ _02730_ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11536__A1 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10339__A2 register_file\[1\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_262_clk clknet_5_19__leaf_clk clknet_leaf_262_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_113_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08952__A2 register_file\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13289__A1 _07660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07982_ _03311_ _03314_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15660__CLK clknet_leaf_135_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09721_ _04894_ register_file\[8\]\[16\] _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11839__A2 _06751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09652_ _04832_ register_file\[23\]\[15\] _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08603_ _03925_ _03929_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09583_ _04893_ _04895_ _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16016__CLK clknet_leaf_229_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15450__A2 register_file\[6\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08534_ _03860_ _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_70_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12264__A2 _07012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13461__A1 _07763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08465_ _03791_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_51_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13213__A1 _07562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08396_ _03723_ _01086_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__A1 _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14961__A1 _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11775__A1 _06266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08640__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13587__I _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09017_ _04336_ _04337_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14713__A1 _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09196__A2 register_file\[24\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15269__A2 register_file\[10\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_253_clk clknet_5_16__leaf_clk clknet_leaf_253_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09919_ _05219_ _05226_ _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15307__I _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11835__I _06718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12930_ _07436_ register_file\[18\]\[19\] _07438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12861_ _07290_ _07391_ _07396_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14600_ _02108_ _01775_ _02109_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11812_ _06741_ register_file\[7\]\[13\] _06742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15580_ _02826_ register_file\[16\]\[23\] _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12792_ _07302_ _07350_ _07354_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16509__CLK clknet_leaf_300_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13452__A1 _07763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10266__A1 _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09120__A2 register_file\[28\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14531_ _02039_ _02041_ _01709_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11743_ _06125_ _06696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14462_ _01058_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12007__A2 register_file\[5\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11674_ _06036_ _06647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16201_ _00589_ clknet_leaf_96_clk register_file\[24\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10018__A1 _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09959__A1 _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13413_ _07734_ register_file\[9\]\[7\] _07741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10625_ _05672_ register_file\[17\]\[30\] _05922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14393_ _01904_ register_file\[30\]\[9\] _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16132_ _00520_ clknet_leaf_76_clk register_file\[31\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13344_ _07534_ _07697_ _07699_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08631__A1 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10556_ _05846_ _05853_ _05854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14704__A1 _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16063_ _00451_ clknet_leaf_306_clk register_file\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10914__I _06169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13275_ _07653_ register_file\[14\]\[16\] _07658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10487_ _05782_ _05785_ _04323_ _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11518__A1 _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15014_ _02518_ register_file\[11\]\[16\] _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15683__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12226_ _06995_ register_file\[31\]\[13\] _06996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14180__A2 register_file\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14830__B _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12191__A1 _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_244_clk clknet_5_17__leaf_clk clknet_leaf_244_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12157_ _06698_ _06943_ _06948_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10741__A2 _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11108_ _06091_ _06286_ _06292_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12088_ _03521_ _06902_ _06906_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16039__CLK clknet_leaf_296_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11039_ _06228_ _06250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15916_ _00304_ clknet_leaf_122_clk register_file\[10\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08698__A1 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12494__A2 _07160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15847_ _00235_ clknet_leaf_46_clk register_file\[12\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15432__A2 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16189__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12246__A2 register_file\[31\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13443__A1 _07553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15778_ _00166_ clknet_leaf_52_clk register_file\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09111__A2 register_file\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14729_ _01986_ register_file\[29\]\[13\] _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08250_ _03576_ _03579_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10009__A1 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08181_ _03274_ register_file\[14\]\[28\] _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08622__A1 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10824__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11509__A1 _06366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10980__A2 _06170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12182__A1 _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_235_clk clknet_5_20__leaf_clk clknet_leaf_235_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08925__A2 register_file\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09834__B _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15120__A1 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07965_ _03051_ register_file\[1\]\[25\] _03052_ _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15127__I register_file\[3\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09704_ _05013_ _05014_ _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08689__A1 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12485__A2 _07153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07896_ _03229_ register_file\[26\]\[25\] _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10496__A1 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09635_ _04945_ _04946_ _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15423__A2 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12237__A2 _07000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09566_ _04877_ _04878_ _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13434__A1 _07543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10248__A1 _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08517_ _03843_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13985__A2 _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09497_ _04810_ register_file\[5\]\[13\] _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11996__A1 _06851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15187__A1 _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08448_ _03768_ _03774_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13737__A2 register_file\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14934__A1 _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08379_ _03706_ register_file\[10\]\[31\] _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_177_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11748__A1 _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10410_ _05710_ _05643_ _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11390_ _06412_ _06472_ _06475_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10341_ _04636_ _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10734__I _06028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10971__A2 register_file\[2\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09169__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13060_ _06048_ _07518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10272_ _05572_ _05573_ _05574_ _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14162__A2 register_file\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12011_ _06815_ register_file\[5\]\[30\] _06860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12173__A1 _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08916__A2 register_file\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_226_clk clknet_5_21__leaf_clk clknet_leaf_226_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_79_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15037__I _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13962_ _01478_ register_file\[30\]\[4\] _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15701_ _00089_ clknet_leaf_211_clk register_file\[28\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12913_ _07422_ register_file\[18\]\[12\] _07428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13893_ _01085_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15414__A2 register_file\[27\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15632_ _00020_ clknet_leaf_165_clk register_file\[30\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12844_ _07274_ _07384_ _07386_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13425__A1 _07742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10239__A1 _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12396__I _07097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15563_ _03060_ _02808_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13976__A2 register_file\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12775_ _07340_ register_file\[20\]\[21\] _07345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16481__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11987__A1 _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14514_ _01161_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11726_ _06103_ _06684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15494_ _01307_ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14925__A1 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14445_ register_file\[5\]\[9\] _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11657_ _06591_ register_file\[10\]\[29\] _06635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11739__A1 _06691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08604__A1 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10608_ _05903_ _05904_ _05905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12400__A2 _07105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14376_ _01880_ _01888_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11588_ _06594_ register_file\[10\]\[0\] _06595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16115_ _00503_ clknet_5_21__leaf_clk register_file\[3\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10411__A1 _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13327_ _07681_ _07689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14116__I _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10539_ _05832_ _05837_ _05838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08080__A2 register_file\[27\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10962__A2 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15350__A1 _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14153__A2 register_file\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16046_ _00434_ clknet_leaf_245_clk register_file\[5\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13258_ _07646_ register_file\[14\]\[9\] _07648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12164__A1 _06706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_217_clk clknet_5_21__leaf_clk clknet_leaf_217_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12209_ _06983_ register_file\[31\]\[8\] _06984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08907__A2 register_file\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09654__B _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13189_ _07538_ _07601_ _07606_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11911__A1 _06796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09580__A2 register_file\[21\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12467__A2 register_file\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10478__A1 _05772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15405__A2 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09420_ _04731_ _04734_ _04529_ _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12219__A2 register_file\[31\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13416__A1 _07742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07894__A2 register_file\[27\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09351_ _03964_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_178_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10819__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11978__A1 _06679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08302_ _01120_ register_file\[27\]\[30\] _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09282_ _04597_ _04598_ _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08233_ _01130_ register_file\[28\]\[29\] _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14916__A1 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10650__A1 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08733__B _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08164_ _03420_ register_file\[23\]\[28\] _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10402__A1 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16204__CLK clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08095_ _03345_ register_file\[9\]\[27\] _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08071__A2 register_file\[23\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10953__A2 _06192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14144__A2 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_208_clk clknet_5_22__leaf_clk clknet_leaf_208_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11902__A1 _06684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input41_I new_value[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16354__CLK clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__A2 register_file\[17\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08997_ _04317_ register_file\[18\]\[6\] _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14447__A3 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ _01178_ _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10469__A1 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07879_ _03213_ _03132_ _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11130__A2 _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07812__B _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09618_ _04661_ register_file\[14\]\[15\] _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10890_ _06155_ _06156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09549_ _04860_ _04861_ _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14080__A1 _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11969__A1 _06830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12560_ _06990_ _07201_ _07203_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__A1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14907__A1 _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10641__A1 _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11511_ _06373_ _06544_ _06548_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12944__I _07417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12491_ _07157_ register_file\[23\]\[16\] _07162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14230_ _01743_ _01488_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14383__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15580__A1 _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11442_ _06382_ _06506_ _06507_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12394__A1 _07102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11197__A2 register_file\[13\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11373_ _06462_ register_file\[26\]\[10\] _06466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14161_ _01110_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08062__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13112_ _06115_ _07555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10324_ _05361_ register_file\[27\]\[25\] _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15332__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14092_ _01147_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12146__A1 _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13043_ _07503_ _07506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10255_ _05359_ register_file\[26\]\[24\] _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13894__A1 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10186_ _05423_ register_file\[13\]\[23\] _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10413__B _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15721__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14994_ _02252_ register_file\[18\]\[16\] _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09314__A2 register_file\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13945_ _01441_ _01462_ _01195_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15399__A1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A2 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13876_ _01146_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15871__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15615_ _00003_ clknet_leaf_19_clk register_file\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12827_ _07257_ _07370_ _07376_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09078__A1 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16595_ _00983_ clknet_leaf_214_clk register_file\[9\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15546_ _03039_ _03044_ _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12758_ _07333_ register_file\[20\]\[14\] _07335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14555__B _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16227__CLK clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11709_ _06081_ _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15477_ _02974_ _02975_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12689_ _07288_ _07284_ _07289_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07948__I _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14428_ _01938_ _01939_ _01859_ _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15571__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11188__A2 register_file\[13\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12385__A1 _07094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14359_ _01871_ _01786_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10935__A2 register_file\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15323__A1 _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14126__A2 register_file\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16377__CLK clknet_leaf_202_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12137__A1 _06933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08920_ _04170_ register_file\[18\]\[5\] _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16029_ _00417_ clknet_leaf_298_clk register_file\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12688__A2 register_file\[21\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13885__A1 _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09553__A2 _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08851_ _04171_ _04173_ _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07802_ _03129_ _03137_ _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08782_ _04031_ register_file\[20\]\[3\] _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09305__A2 _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_4__f_clk clknet_3_1_0_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_22_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11112__A2 register_file\[27\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12860__A2 register_file\[1\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09403_ _04714_ _04717_ _04018_ _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10871__A1 _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14062__A1 _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09334_ _04582_ register_file\[4\]\[11\] _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08019__I _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09265_ _03863_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08292__A2 register_file\[22\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08216_ _01081_ register_file\[20\]\[29\] _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09196_ _04239_ register_file\[24\]\[9\] _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11179__A2 _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12376__A1 _07090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08147_ _03320_ register_file\[31\]\[28\] _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09241__A1 _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10926__A2 _06178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08078_ _03409_ _03163_ _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12128__A1 _06670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15744__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12679__A2 _07272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10040_ _05342_ _05345_ _04675_ _05346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11351__A2 _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12939__I _07406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11991_ _06844_ register_file\[5\]\[21\] _06849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11103__A2 _06286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12300__A1 _06969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13730_ _01249_ register_file\[10\]\[1\] _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10942_ _06189_ register_file\[2\]\[14\] _06191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07858__A2 _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12851__A2 _07384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09313__I _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13661_ _01179_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10873_ net29 _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15400_ _02818_ register_file\[21\]\[21\] _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12612_ _07234_ _07235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16380_ _00768_ clknet_leaf_278_clk register_file\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12603__A2 register_file\[22\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13592_ _01109_ _01112_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15331_ _02581_ register_file\[19\]\[20\] _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10614__A1 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12543_ _07185_ _07193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12674__I _07231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09480__A1 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08283__A2 _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15262_ _01079_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12474_ _07150_ register_file\[23\]\[9\] _07152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12367__A1 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14213_ _01726_ _01468_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11425_ _06495_ _06496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09232__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15193_ _02694_ _02609_ _02695_ _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08035__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10917__A2 register_file\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15305__A1 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14144_ _01658_ _01490_ _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14108__A2 register_file\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09783__A2 register_file\[30\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11356_ _06377_ _06448_ _06455_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07794__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10307_ _03907_ _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_193_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14075_ _01508_ register_file\[8\]\[5\] _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11287_ _06094_ _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13026_ _07295_ _07494_ _07495_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10238_ _05539_ _05540_ _05541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11342__A2 _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15608__A2 register_file\[11\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10169_ _05340_ register_file\[24\]\[23\] _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13619__A1 _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09299__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14977_ _02480_ _02481_ _02399_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11753__I _06138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13928_ register_file\[4\]\[3\] _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12842__A2 _07384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13859_ _01202_ register_file\[16\]\[3\] _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15617__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16578_ _00966_ clknet_leaf_14_clk register_file\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15529_ _03027_ register_file\[13\]\[22\] _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09050_ _04369_ register_file\[12\]\[7\] _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12358__A1 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08001_ _03003_ register_file\[28\]\[26\] _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15767__CLK clknet_leaf_224_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09223__A1 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08026__A2 _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11030__A1 _06240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09952_ _05257_ _05258_ _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10832__I _06025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13858__A1 _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08903_ _04225_ _03929_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09883_ _05190_ register_file\[26\]\[19\] _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11333__A2 _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08834_ _04157_ _03929_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08765_ _04087_ _04088_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_263_clk_I clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13086__A2 register_file\[16\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11663__I _06020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12833__A2 register_file\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08696_ _03803_ register_file\[20\]\[2\] _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10844__A1 _06109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14035__A1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08972__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_278_clk_I clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16542__CLK clknet_leaf_302_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12597__A1 _07219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09317_ _04633_ register_file\[1\]\[10\] _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14338__A2 register_file\[9\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09248_ _04499_ register_file\[3\]\[9\] _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_201_clk_I clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12349__A1 _07018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09214__A1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09179_ _04288_ register_file\[2\]\[8\] _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13010__A2 register_file\[17\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11021__A1 _06082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11210_ _06126_ _06351_ _06354_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12190_ _06962_ _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07776__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11572__A2 _06582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10742__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11141_ _06152_ _06307_ _06311_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput44 net44 rD[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_clkbuf_leaf_216_clk_I clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput55 net55 rD[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__13849__A1 _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output72_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput66 net66 rD[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09517__A2 register_file\[10\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput77 net77 rS[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11072_ _06270_ _06271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_110_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput88 net88 rS[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_62_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput99 net99 rS[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_66_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12521__A1 _07135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11324__A2 _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14900_ _02321_ register_file\[30\]\[15\] _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10023_ _05061_ register_file\[5\]\[21\] _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15880_ _00268_ clknet_leaf_109_clk register_file\[11\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14831_ _02333_ _02337_ _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13077__A2 _07520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11088__A1 _06275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14762_ _01423_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11974_ _06837_ register_file\[5\]\[14\] _06839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12824__A2 register_file\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16501_ _00889_ clknet_leaf_225_clk register_file\[15\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13713_ _01231_ _01084_ _01232_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14884__I _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10925_ _06174_ register_file\[2\]\[7\] _06181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14693_ register_file\[7\]\[12\] _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14026__A1 _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16432_ _00820_ clknet_leaf_161_clk register_file\[17\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13644_ register_file\[5\]\[0\] _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14577__A2 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10856_ net26 _06128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12588__A1 _07219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16363_ _00751_ clknet_leaf_140_clk register_file\[1\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09453__A1 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13575_ _01095_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08256__A2 _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10787_ _06071_ _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15314_ _02811_ _02813_ _02814_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14329__A2 register_file\[21\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15526__A1 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12526_ _07036_ _07138_ _07181_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16294_ _00682_ clknet_leaf_80_clk register_file\[21\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15245_ _02745_ _02746_ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12457_ _06967_ _07136_ _07141_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09205__A1 _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13001__A2 register_file\[17\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11012__A1 _06064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11408_ _06457_ _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09756__A2 register_file\[18\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15176_ _02675_ _02678_ _02508_ _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12388_ _06978_ _07098_ _07100_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14127_ _01557_ register_file\[26\]\[6\] _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11339_ _06442_ _06371_ _06443_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09508__A2 register_file\[30\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14058_ _01308_ register_file\[17\]\[5\] _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13963__I _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13009_ _07278_ _07480_ _07485_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16415__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14265__A1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11483__I _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08550_ _03876_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16565__CLK clknet_leaf_215_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08481_ _03807_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09692__A1 _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12579__A1 _07009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09444__A1 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13240__A2 register_file\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09102_ _04418_ _04421_ _03961_ _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11251__A1 _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15517__A1 _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09033_ _04213_ register_file\[12\]\[6\] _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09747__A2 register_file\[27\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14740__A2 _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12751__A1 _07326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14034__I _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09935_ _05227_ _05242_ _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14969__I _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16095__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12503__A1 _07164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09866_ _04970_ register_file\[1\]\[18\] _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08817_ _04132_ _04140_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09797_ _04970_ register_file\[1\]\[17\] _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14256__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13059__A2 _07505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_82_clk_I clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ _04071_ _04072_ _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12806__A2 register_file\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10817__A1 _06087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09683__A1 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08679_ _03920_ register_file\[3\]\[1\] _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10710_ _03883_ register_file\[12\]\[31\] _06006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14559__A2 _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11490__A1 _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11690_ _06650_ register_file\[8\]\[6\] _06659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_97_clk_I clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10641_ _05756_ register_file\[21\]\[30\] _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10737__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08238__A2 _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_140_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13113__I _07519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13231__A2 _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13360_ _07708_ register_file\[29\]\[18\] _07709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10572_ _05854_ _05869_ _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07997__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12311_ _07041_ _07054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12990__A1 _07259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_20_clk_I clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11793__A2 register_file\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13291_ _07630_ _07667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15030_ register_file\[7\]\[16\] _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12242_ _06959_ _07007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14731__A2 register_file\[30\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_155_clk_I clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11568__I _06553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12742__A1 _07252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16438__CLK clknet_leaf_204_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12173_ _06911_ register_file\[3\]\[31\] _06957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_35_clk_I clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11124_ _06297_ register_file\[27\]\[21\] _06302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13298__A2 _07670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15932_ _00320_ clknet_leaf_287_clk register_file\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11055_ _06144_ _06257_ _06259_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08174__A1 _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16588__CLK clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10006_ _03934_ _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15863_ _00251_ clknet_leaf_223_clk register_file\[12\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14814_ _01071_ _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15794_ _00182_ clknet_leaf_168_clk register_file\[19\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14745_ _02252_ register_file\[18\]\[13\] _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11957_ _06822_ register_file\[5\]\[7\] _06829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09674__A1 _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13470__A2 _07730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11481__A1 _06524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10908_ _06170_ register_file\[2\]\[0\] _06171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14676_ _02184_ _01853_ _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11888_ _06670_ _06785_ _06787_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16415_ _00803_ clknet_leaf_15_clk register_file\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13627_ _01147_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10839_ _06113_ _06096_ _06114_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_108_clk_I clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08229__A2 register_file\[27\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13222__A2 _07622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16346_ _00734_ clknet_leaf_270_clk register_file\[20\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13558_ _00992_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09977__A2 register_file\[6\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14970__A2 register_file\[24\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07988__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13958__I _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12981__A1 _07462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12509_ _07018_ _07167_ _07172_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16277_ _00665_ clknet_leaf_208_clk register_file\[22\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13489_ _01009_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15228_ _02728_ _02729_ _02399_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11536__A2 _06561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12733__A1 _07318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15159_ _02576_ register_file\[25\]\[18\] _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15278__A3 _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15805__CLK clknet_leaf_279_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07981_ _03312_ _03313_ _03231_ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13289__A2 register_file\[14\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09720_ _04892_ register_file\[9\]\[16\] _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09651_ _04830_ register_file\[22\]\[15\] _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14238__A1 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15955__CLK clknet_leaf_226_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08602_ _03928_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09582_ _04894_ register_file\[20\]\[14\] _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14789__A2 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08533_ _03798_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13461__A2 register_file\[9\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11472__A1 _06524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08464_ net4 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15202__A3 _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09417__A1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13213__A2 _07615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08395_ register_file\[31\]\[31\] _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14410__A1 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11224__A1 _06152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10027__A2 register_file\[6\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14961__A2 register_file\[1\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07979__A1 _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11775__A2 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12972__A1 _07241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12772__I _07321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09016_ _04125_ register_file\[8\]\[6\] _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12724__A1 _07314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14699__I register_file\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09918_ _05222_ _05225_ _03992_ _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08156__A1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09849_ _05023_ register_file\[18\]\[18\] _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12860_ _07395_ register_file\[1\]\[23\] _07396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11811_ _06721_ _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09656__A1 _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12791_ _07311_ register_file\[20\]\[28\] _07354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13452__A2 register_file\[9\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14530_ _02040_ _01707_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11463__A1 _06405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10266__A2 register_file\[31\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11742_ _06694_ _06692_ _06695_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14461_ _01635_ register_file\[24\]\[10\] _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09408__A1 _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11673_ _06645_ _06641_ _06646_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16200_ _00588_ clknet_leaf_92_clk register_file\[24\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10018__A2 register_file\[18\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11215__A1 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13412_ _07522_ _07738_ _07740_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10624_ _05917_ _05920_ _04183_ _05921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14392_ _01071_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14952__A2 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16131_ _00519_ clknet_leaf_61_clk register_file\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13343_ _07694_ register_file\[29\]\[11\] _07699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16260__CLK clknet_leaf_75_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10555_ _05849_ _05852_ _03856_ _05853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16062_ _00450_ clknet_leaf_300_clk register_file\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15828__CLK clknet_leaf_172_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13274_ _07543_ _07656_ _07657_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14704__A2 register_file\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10486_ _05783_ _05784_ _05785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11298__I _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15013_ _01681_ _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12715__A1 _07306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11518__A2 _06544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12225_ _06962_ _06995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12191__A2 register_file\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12156_ _06947_ register_file\[3\]\[23\] _06948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14468__A1 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11107_ _06290_ register_file\[27\]\[14\] _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15978__CLK clknet_leaf_291_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14402__I _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12087_ _06863_ net31 _06906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08147__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13140__A1 _07504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11038_ _06113_ _06243_ _06249_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15915_ _00303_ clknet_leaf_112_clk register_file\[10\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08698__A2 register_file\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15846_ _00234_ clknet_leaf_47_clk register_file\[12\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09647__A1 _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12989_ _07470_ register_file\[17\]\[10\] _07474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15777_ _00165_ clknet_leaf_52_clk register_file\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13443__A2 _07752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11454__A1 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14728_ _02235_ register_file\[28\]\[13\] _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14659_ _02163_ _02167_ _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15196__A2 _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_180_clk clknet_5_29__leaf_clk clknet_leaf_180_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_177_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16603__CLK clknet_leaf_284_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10009__A2 register_file\[20\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11206__A1 _06117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08180_ _03509_ _03436_ _03510_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14293__B _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12954__A1 _07304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12592__I _07193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16329_ _00717_ clknet_leaf_99_clk register_file\[20\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08622__A2 register_file\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10326__B _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12706__A1 _07300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11509__A2 _06544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08386__A1 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12182__A2 _06961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10193__A1 _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11936__I _06814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14312__I _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ _03294_ _03295_ _03297_ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_190_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09703_ _04812_ register_file\[16\]\[16\] _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13131__A1 _07563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07895_ _01042_ _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09634_ _04812_ register_file\[4\]\[15\] _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10496__A2 register_file\[5\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11693__A1 _06650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16133__CLK clknet_leaf_79_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12767__I _07310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09565_ _04812_ register_file\[8\]\[14\] _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15143__I _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14631__A1 _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13434__A2 _07752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11671__I _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11445__A1 _06502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08516_ _03770_ _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10248__A2 register_file\[6\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09496_ _03840_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_169_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08310__A1 _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08447_ _03773_ register_file\[24\]\[0\] _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10287__I _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_171_clk clknet_5_28__leaf_clk clknet_leaf_171_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__15187__A2 register_file\[10\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13198__A1 _07548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14934__A2 register_file\[13\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08378_ _01277_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_177_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13598__I _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11748__A2 register_file\[8\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12945__A1 _07443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09297__B _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09810__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10340_ _05638_ _05639_ _05641_ _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14931__B _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14698__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10271_ _05306_ register_file\[1\]\[24\] _05574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13370__A1 _07560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12010_ _06712_ _06854_ _06859_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12173__A2 register_file\[3\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10750__I _06028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15111__A2 _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09316__I _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13961_ _01042_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12912_ _07262_ _07425_ _07427_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15700_ _00088_ clknet_leaf_179_clk register_file\[28\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13892_ _01083_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14378__B _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12843_ _07381_ register_file\[1\]\[16\] _07386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12677__I _06112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15631_ _00019_ clknet_leaf_152_clk register_file\[30\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14622__A1 _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15562_ _03058_ _03059_ _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10239__A2 register_file\[14\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11436__A1 _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12774_ _07283_ _07343_ _07344_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14513_ _02022_ _01775_ _02023_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11987__A2 _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11725_ _06682_ _06680_ _06683_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10197__I _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15493_ _02826_ register_file\[24\]\[22\] _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_162_clk clknet_5_31__leaf_clk clknet_leaf_162_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13189__A1 _07538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08890__I _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14444_ _01954_ _01955_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14925__A2 register_file\[9\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11656_ _06438_ _06630_ _06634_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15650__CLK clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12936__A1 _07286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11739__A2 _06692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10607_ _03920_ register_file\[11\]\[30\] _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14375_ _01887_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11587_ _06593_ _06594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_128_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16114_ _00502_ clknet_leaf_229_clk register_file\[3\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13326_ _07516_ _07680_ _07688_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_182_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10538_ _05836_ _05643_ _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__16006__CLK clknet_leaf_309_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16045_ _00433_ clknet_leaf_249_clk register_file\[5\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13257_ _07526_ _07642_ _07647_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10469_ _05501_ register_file\[26\]\[27\] _05769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08368__A1 _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12208_ _06962_ _06983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13361__A1 _07550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12164__A2 _06950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13188_ _07605_ register_file\[15\]\[13\] _07606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10175__A1 _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11911__A2 register_file\[6\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12139_ _06933_ register_file\[3\]\[16\] _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16156__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13971__I _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11675__A1 _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14288__B _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12587__I _07182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15829_ _00217_ clknet_leaf_219_clk register_file\[26\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13416__A2 register_file\[9\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14613__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09350_ _04660_ _04665_ _03838_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08301_ _03629_ _01117_ _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11978__A2 _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09281_ _04327_ register_file\[16\]\[10\] _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_153_clk clknet_5_30__leaf_clk clknet_leaf_153_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_166_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08232_ _03558_ _03561_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14916__A2 register_file\[21\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10835__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08163_ _01123_ register_file\[22\]\[28\] _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13211__I _07582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08094_ _03181_ register_file\[8\]\[27\] _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09845__B _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08359__A1 _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_19__f_clk_I clknet_3_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11666__I _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11902__A2 _06792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08996_ _04316_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13104__A1 _07548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input34_I new_value[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08040__I register_file\[5\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07947_ _03270_ _03280_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14852__A1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10469__A2 register_file\[26\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07878_ register_file\[3\]\[24\] _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09617_ _04927_ _04928_ _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07885__A3 _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11418__A1 _06440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09548_ _04729_ register_file\[28\]\[14\] _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15673__CLK clknet_leaf_241_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11969__A2 register_file\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12091__A1 _06863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_144_clk clknet_5_27__leaf_clk clknet_leaf_144_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09479_ _04785_ _04792_ _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08834__A2 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11510_ _06546_ register_file\[11\]\[1\] _06548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12490_ _06999_ _07160_ _07161_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14907__A2 register_file\[17\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10641__A2 register_file\[21\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12918__A1 _07429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11441_ _06502_ register_file\[12\]\[5\] _06507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15580__A2 register_file\[16\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12394__A2 register_file\[24\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13591__A1 _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14160_ _01508_ register_file\[8\]\[6\] _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11372_ _06457_ _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_180_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13111_ _07553_ _07544_ _07554_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10323_ _05359_ register_file\[26\]\[25\] _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12960__I _07454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14091_ _01604_ _01258_ _01606_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15332__A2 register_file\[18\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16179__CLK clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13343__A1 _07694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13042_ _07504_ _07505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10254_ _05555_ _05556_ _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10157__A1 _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13894__A2 register_file\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10185_ _05485_ _05488_ _05421_ _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15096__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14887__I _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14993_ _02164_ register_file\[19\]\[16\] _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14843__A1 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11657__A1 _06591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13944_ _01452_ _01461_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15399__A2 register_file\[20\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13875_ _01391_ _01046_ _01392_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_165_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12826_ _07374_ register_file\[1\]\[9\] _07376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15614_ _00002_ clknet_leaf_24_clk register_file\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11409__A1 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16594_ _00982_ clknet_leaf_176_clk register_file\[9\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14071__A2 _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12757_ _07266_ _07329_ _07334_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15545_ _03041_ _03043_ _02960_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_135_clk clknet_5_26__leaf_clk clknet_leaf_135_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15511__I _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11708_ _06670_ _06668_ _06671_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15476_ _02805_ register_file\[17\]\[22\] _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12688_ _07279_ register_file\[21\]\[22\] _07289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15020__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12909__A1 _07422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14427_ _01684_ register_file\[10\]\[9\] _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11639_ _06620_ register_file\[10\]\[21\] _06625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15571__A2 register_file\[28\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12385__A2 register_file\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14358_ register_file\[7\]\[8\] _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_183_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13309_ _07631_ register_file\[14\]\[31\] _07677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14289_ _01799_ _01802_ _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13334__A1 _07524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16028_ _00416_ clknet_leaf_293_clk register_file\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13885__A2 register_file\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08850_ _04172_ register_file\[19\]\[4\] _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15087__A1 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07801_ _03136_ _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08781_ _04029_ register_file\[21\]\[3\] _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15696__CLK clknet_leaf_165_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10320__A1 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07867__A3 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09402_ _04715_ _04716_ _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10871__A2 register_file\[30\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14746__B _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09333_ _04580_ register_file\[5\]\[11\] _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12073__A1 _06892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_126_clk clknet_5_25__leaf_clk clknet_leaf_126_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_34_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08744__B _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09264_ _04580_ register_file\[21\]\[10\] _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11820__A1 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08215_ _03541_ _03544_ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14037__I _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09195_ _04237_ register_file\[25\]\[9\] _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14365__A3 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08146_ _03153_ register_file\[30\]\[28\] _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16321__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09241__A2 register_file\[28\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08044__A3 _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13876__I _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14117__A3 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08077_ _03407_ _03408_ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12128__A2 _06929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13325__A1 _07686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11396__I _06457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16471__CLK clknet_leaf_215_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11887__A1 _06782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15078__A1 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08979_ _01706_ _03763_ _04299_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11639__A1 _06620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11990_ _06691_ _06847_ _06848_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12300__A2 _07040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10941_ _06086_ _06185_ _06190_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13116__I _06120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13660_ register_file\[3\]\[0\] _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10872_ _06139_ _06140_ _06141_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14053__A2 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12611_ _07231_ _07234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12064__A1 _06892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_117_clk clknet_5_24__leaf_clk clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13591_ _01111_ register_file\[9\]\[0\] _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15330_ _02830_ _01010_ _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12542_ _06972_ _07184_ _07192_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09480__A2 register_file\[17\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15261_ _02742_ _02761_ _02762_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12473_ _06982_ _07146_ _07151_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14212_ _01725_ _01553_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11424_ _06494_ _06495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_184_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15192_ _02610_ register_file\[13\]\[18\] _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09232__A2 register_file\[18\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14143_ _01657_ _01488_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12690__I _06129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11355_ _06454_ register_file\[26\]\[3\] _06455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15305__A2 register_file\[25\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13316__A1 _07682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08991__A1 _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10306_ _05607_ register_file\[14\]\[25\] _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07794__A2 register_file\[2\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14074_ _01571_ _01589_ _01506_ _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11286_ _06405_ _06396_ _06406_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13025_ _07491_ register_file\[17\]\[25\] _07495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10237_ _05340_ register_file\[12\]\[24\] _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11878__A1 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10168_ _05338_ register_file\[25\]\[23\] _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13619__A2 register_file\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10550__A1 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10099_ _05338_ register_file\[21\]\[22\] _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09299__A2 register_file\[24\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14976_ _02397_ register_file\[26\]\[16\] _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13927_ _01442_ _01444_ _01266_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10302__A1 _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13858_ _01332_ _01376_ _01201_ net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15241__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12809_ _07239_ _07360_ _07365_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_108_clk clknet_5_12__leaf_clk clknet_leaf_108_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16577_ _00965_ clknet_leaf_14_clk register_file\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13789_ _01307_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15528_ _01047_ _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11802__A1 _06734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16344__CLK clknet_leaf_195_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12086__B _06905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15459_ _02957_ _02958_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08000_ _03329_ _03332_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12358__A2 _07078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15397__B _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09223__A2 register_file\[8\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13696__I _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16494__CLK clknet_leaf_188_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13307__A1 _07631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07785__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09951_ _05192_ register_file\[19\]\[20\] _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10334__B _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08902_ _04222_ _04223_ _04224_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09882_ _03807_ _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08833_ _04153_ _04155_ _04156_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14807__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08764_ _03773_ register_file\[12\]\[3\] _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09414__I _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12294__A1 _07042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08695_ _03800_ register_file\[21\]\[2\] _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10844__A2 register_file\[30\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15232__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14035__A2 register_file\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07869__I register_file\[4\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09316_ _03922_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10509__B _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09247_ _04288_ register_file\[2\]\[9\] _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15711__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12349__A2 _07071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _04491_ _04496_ _04220_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09214__A2 register_file\[20\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ _03458_ _03460_ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11021__A2 _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07776__A2 register_file\[13\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08973__A1 _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11140_ _06268_ register_file\[27\]\[28\] _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10780__A1 _06064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput45 net45 rD[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput56 net56 rD[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput67 net67 rD[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_27_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11071_ _06267_ _06270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput78 net78 rS[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_89_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput89 net89 rS[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output65_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08725__A1 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10022_ _05320_ _05327_ _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12521__A2 register_file\[23\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16217__CLK clknet_leaf_196_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14830_ _02334_ _02335_ _02336_ _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09324__I _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14761_ _02267_ _02268_ _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11088__A2 register_file\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12285__A1 _06960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11973_ _06674_ _06833_ _06838_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09150__A1 _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16500_ _00888_ clknet_leaf_174_clk register_file\[15\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10924_ _06056_ _06178_ _06180_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13712_ _01086_ register_file\[29\]\[1\] _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14692_ _02033_ register_file\[6\]\[12\] _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_45_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16367__CLK clknet_leaf_144_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14386__B _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16431_ _00819_ clknet_leaf_144_clk register_file\[17\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12037__A1 _06870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10855_ _06126_ _06118_ _06127_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13643_ _01162_ _01163_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08384__B _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16362_ _00750_ clknet_leaf_96_clk register_file\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13574_ _00997_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10786_ net12 _06071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09453__A2 register_file\[15\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15313_ _01559_ _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12525_ _07135_ register_file\[23\]\[31\] _07181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16293_ _00681_ clknet_leaf_75_clk register_file\[21\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15526__A2 register_file\[12\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15244_ _01114_ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12456_ _07138_ register_file\[23\]\[2\] _07141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08008__A3 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09205__A2 register_file\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11407_ _06429_ _06479_ _06485_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11012__A2 _06229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15175_ _02676_ _02592_ _02677_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12387_ _07094_ register_file\[24\]\[6\] _07100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14126_ _01382_ register_file\[27\]\[6\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11338_ _06368_ register_file\[19\]\[30\] _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14057_ _01572_ register_file\[16\]\[5\] _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11269_ _06393_ _06384_ _06394_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14501__A3 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13008_ _07484_ register_file\[17\]\[18\] _07485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10523__A1 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15236__I _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14265__A2 register_file\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12276__A1 _06960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14959_ _02464_ _02300_ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08480_ _03806_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_78_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15214__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12579__A2 _07208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13776__A1 _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09101_ _04419_ _04420_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15517__A2 register_file\[8\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11251__A2 _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09032_ _04211_ register_file\[13\]\[6\] _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13528__A1 _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11939__I _06817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10843__I _06051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12200__A1 _06974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08955__A1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12751__A2 register_file\[20\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09934_ _05236_ _05241_ _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08707__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12503__A2 register_file\[23\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09865_ _05173_ register_file\[3\]\[18\] _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11674__I _06036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09380__A1 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08183__A2 _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08816_ _04135_ _04138_ _04139_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09796_ _04837_ register_file\[3\]\[17\] _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12267__A1 _07019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08747_ _03901_ register_file\[28\]\[2\] _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ _03917_ register_file\[2\]\[1\] _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output103_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11490__A2 _06534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10640_ _05933_ _05936_ _03914_ _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10571_ _05861_ _05868_ _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12310_ _06980_ _07050_ _07053_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13519__A1 _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07997__A2 register_file\[27\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12990__A2 _07473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13290_ _07560_ _07663_ _07666_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09199__A1 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12241_ _06107_ _07006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10753__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__I _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12742__A2 _07322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12172_ _06714_ _06914_ _06956_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08410__A3 _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11123_ _06117_ _06300_ _06301_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14495__A2 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11054_ _06254_ register_file\[28\]\[26\] _06259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15931_ _00319_ clknet_leaf_265_clk register_file\[10\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11584__I _06590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09371__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10005_ _05295_ _05311_ _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_188_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15862_ _00250_ clknet_leaf_220_clk register_file\[12\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15444__A1 _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07921__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14813_ _02317_ _02318_ _02319_ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15793_ _00181_ clknet_leaf_168_clk register_file\[19\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15757__CLK clknet_leaf_148_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09123__A1 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14744_ _01404_ _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11956_ _06658_ _06826_ _06828_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_189_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09674__A2 register_file\[21\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10907_ _06169_ _06170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_162_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11481__A2 register_file\[12\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14675_ _02182_ _02183_ _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11887_ _06782_ register_file\[6\]\[11\] _06787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16414_ _00802_ clknet_leaf_27_clk register_file\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10838_ _06109_ register_file\[30\]\[19\] _06114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09003__B _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13626_ _01146_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12430__A1 _07123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16345_ _00733_ clknet_leaf_196_clk register_file\[20\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10769_ _06056_ _06052_ _06057_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13557_ _01067_ _01077_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07988__A2 register_file\[23\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12981__A2 register_file\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12508_ _07171_ register_file\[23\]\[23\] _07172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13488_ _01008_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16276_ _00664_ clknet_leaf_208_clk register_file\[22\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10992__A1 _06021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_262_clk_I clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14135__I _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15227_ _02397_ register_file\[18\]\[19\] _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12439_ _07087_ register_file\[24\]\[28\] _07130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12733__A2 register_file\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15158_ _02411_ register_file\[24\]\[18\] _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08401__A3 _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14109_ register_file\[3\]\[5\] _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15089_ _01142_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09673__B _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07980_ _03229_ register_file\[18\]\[26\] _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_277_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16532__CLK clknet_leaf_174_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12497__A1 _07006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08165__A2 _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09650_ _04960_ _04961_ _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14238__A2 register_file\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15435__A1 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08601_ _03927_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_110_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09581_ _03882_ _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08532_ _03819_ _03858_ _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13997__A1 _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08463_ _03789_ _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_215_clk_I clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13749__A1 _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08394_ _03701_ register_file\[30\]\[31\] _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_177_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14410__A2 register_file\[20\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12421__A1 _07116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11224__A2 _06358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_clk clknet_5_6__leaf_clk clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_177_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12972__A2 _07456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09015_ _04122_ register_file\[9\]\[6\] _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14174__A1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16062__CLK clknet_leaf_300_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08928__A1 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08043__I _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10735__A1 _06029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14477__A2 _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09917_ _05223_ _05224_ _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_97_clk clknet_5_15__leaf_clk clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08156__A2 register_file\[19\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09848_ _05155_ _05156_ _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11160__A1 _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07903__A2 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09779_ _05088_ register_file\[29\]\[17\] _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09105__A1 _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15604__I _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11810_ _06672_ _06737_ _06740_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12790_ _07300_ _07350_ _07353_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09656__A2 register_file\[2\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11741_ _06687_ register_file\[8\]\[21\] _06695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11463__A2 _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14460_ _01931_ _01971_ _01634_ net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11672_ _06643_ register_file\[8\]\[1\] _06646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09408__A2 register_file\[31\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13411_ _07734_ register_file\[9\]\[6\] _07740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10623_ _05918_ _05919_ _05920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12412__A1 _07002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14391_ _01900_ _01901_ _01902_ _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11215__A2 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12963__I _07457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16405__CLK clknet_leaf_213_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13342_ _07531_ _07697_ _07698_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16130_ _00518_ clknet_leaf_60_clk register_file\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10554_ _05850_ _05851_ _05852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10974__A1 _06148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13273_ _07653_ register_file\[14\]\[15\] _07657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16061_ _00449_ clknet_leaf_300_clk register_file\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10485_ _05583_ register_file\[19\]\[28\] _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09049__I _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12224_ _06085_ _06994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15012_ _02516_ _02272_ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12715__A2 _07235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13912__A1 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13794__I _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09493__B _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12155_ _06910_ _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08888__I _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14468__A2 register_file\[27\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11106_ _06086_ _06286_ _06291_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12479__A1 _07150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12086_ _03448_ _06902_ _06905_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_88_clk clknet_5_14__leaf_clk clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08147__A2 register_file\[31\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11037_ _06247_ register_file\[28\]\[19\] _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15914_ _00302_ clknet_leaf_112_clk register_file\[10\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13140__A2 register_file\[16\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11151__A1 _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15845_ _00233_ clknet_leaf_61_clk register_file\[12\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__B _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15776_ _00164_ clknet_leaf_13_clk register_file\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12988_ _07465_ _07473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09647__A2 _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14727_ _01080_ _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12651__A1 _07255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11454__A2 _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11939_ _06817_ _06818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14658_ _02165_ _02166_ _01919_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11206__A2 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13609_ _01129_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16085__CLK clknet_leaf_233_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14589_ _02098_ _01853_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_12_clk clknet_5_2__leaf_clk clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16328_ _00716_ clknet_leaf_79_clk register_file\[20\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12954__A2 _07446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10965__A1 _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_81_clk_I clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16259_ _00647_ clknet_leaf_78_clk register_file\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12706__A2 _07296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13903__A1 _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10717__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08798__I _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11390__A1 _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10193__A2 _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_96_clk_I clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07963_ _03296_ _03132_ _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_79_clk clknet_5_11__leaf_clk clknet_leaf_79_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08138__A2 _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09702_ _04810_ register_file\[17\]\[16\] _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13131__A2 register_file\[16\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07894_ _03063_ register_file\[27\]\[25\] _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15408__A1 _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11142__A1 _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09633_ _04810_ register_file\[5\]\[15\] _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11693__A2 register_file\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15424__I _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11952__I _06825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09564_ _04810_ register_file\[9\]\[14\] _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_1__f_clk_I clknet_3_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_154_clk_I clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08515_ _03841_ register_file\[17\]\[0\] _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12642__A1 _07254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09495_ _04793_ _04808_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16428__CLK clknet_leaf_140_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08310__A2 register_file\[31\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_clk_I clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08446_ _03772_ _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08038__I register_file\[4\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14395__A1 _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13198__A2 _07608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08377_ _03702_ _03704_ _01170_ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_169_clk_I clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12945__A2 register_file\[18\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16578__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09810__A2 register_file\[23\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_49_clk_I clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07821__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10270_ _05508_ register_file\[3\]\[24\] _05573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10708__A1 _05996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09574__A1 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13370__A2 _07711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11381__A1 _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08501__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09326__A1 _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_107_clk_I clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13119__I _06124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13960_ _01474_ _01475_ _01476_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_150_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12911_ _07422_ register_file\[18\]\[11\] _07427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13891_ _01319_ register_file\[28\]\[3\] _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15630_ _00018_ clknet_leaf_152_clk register_file\[30\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12842_ _07271_ _07384_ _07385_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14622__A2 register_file\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15561_ _02805_ register_file\[25\]\[23\] _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11436__A2 _06496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12773_ _07340_ register_file\[20\]\[20\] _07344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08301__A2 _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14512_ _01776_ register_file\[13\]\[10\] _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11724_ _06675_ register_file\[8\]\[16\] _06683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15492_ _02983_ _02990_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15178__A3 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13789__I _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13189__A2 _07601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14443_ register_file\[4\]\[9\] _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11655_ _06591_ register_file\[10\]\[28\] _06634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08392__B _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12936__A2 _07439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10606_ _03828_ register_file\[10\]\[30\] _05903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14374_ _01885_ _01886_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11586_ _06590_ _06593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10947__A1 _06189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10427__B _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16113_ _00501_ clknet_leaf_226_clk register_file\[3\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10537_ _05833_ _05834_ _05835_ _05836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_13325_ _07686_ register_file\[29\]\[4\] _07688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15945__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14689__A2 _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16044_ _00432_ clknet_leaf_251_clk register_file\[5\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13256_ _07646_ register_file\[14\]\[8\] _07647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10468_ _05766_ _05767_ _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09565__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12207_ _06063_ _06982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13361__A2 _07704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13187_ _07585_ _07605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10399_ _05563_ register_file\[9\]\[26\] _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10175__A2 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12138_ _06679_ _06936_ _06937_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_170_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__A1 _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14310__A1 _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12069_ _06892_ net23 _06896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11124__A1 _06297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_1_clk clknet_5_0__leaf_clk clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09868__A2 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11675__A2 register_file\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12872__A1 _07302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11772__I _06163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15244__I _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15828_ _00216_ clknet_leaf_172_clk register_file\[26\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15759_ _00147_ clknet_leaf_146_clk register_file\[13\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12624__A1 _07241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08300_ _03628_ _01115_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09280_ _04325_ register_file\[17\]\[10\] _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08231_ _03559_ _03560_ _01126_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08162_ _03491_ _01133_ _03492_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10938__A1 _06082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07803__A1 _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08093_ _03406_ _03424_ _03179_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_146_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15341__A3 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11363__A1 _06454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16100__CLK clknet_leaf_54_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08995_ _03778_ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14301__A1 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13104__A2 _07544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07946_ _03273_ _03278_ _03279_ _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11115__A1 _06104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input27_I new_value[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12863__A1 _07293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ _02964_ register_file\[2\]\[24\] _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_99_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16250__CLK clknet_leaf_269_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09616_ _04729_ register_file\[12\]\[15\] _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14604__A2 _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09152__I _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09547_ _04727_ register_file\[29\]\[14\] _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11418__A2 _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08295__A1 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09478_ _04788_ _04791_ _04382_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12091__A2 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14368__A1 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08429_ _03754_ _03756_ _01170_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15968__CLK clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13402__I _07729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12918__A2 register_file\[18\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11440_ _06505_ _06506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13040__A1 _06216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10929__A1 _06064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09795__A1 _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11371_ _06393_ _06458_ _06464_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12018__I _06862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output95_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13110_ _07551_ register_file\[16\]\[19\] _07554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10322_ _05622_ _05623_ _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14090_ _01605_ register_file\[15\]\[5\] _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11857__I _06767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09547__A1 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13041_ _07503_ _07504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10761__I _06028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13343__A2 register_file\[29\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10253_ _05425_ register_file\[24\]\[24\] _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_29__f_clk clknet_3_7_0_clk clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10157__A2 register_file\[19\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10184_ _05486_ _05487_ _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11106__A1 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14992_ _02496_ _02249_ _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14843__A2 register_file\[8\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13943_ _01460_ _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12854__A1 _07283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13874_ _01216_ register_file\[23\]\[3\] _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09062__I _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15613_ _00001_ clknet_leaf_32_clk register_file\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12825_ _07254_ _07370_ _07375_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12606__A1 _07036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11409__A2 register_file\[26\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16593_ _00981_ clknet_leaf_178_clk register_file\[9\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15544_ _03042_ _02958_ _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08286__A1 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12756_ _07333_ register_file\[20\]\[13\] _07334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12082__A2 _06902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10093__A1 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11707_ _06663_ register_file\[8\]\[11\] _06671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15475_ _02889_ register_file\[16\]\[22\] _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12687_ _06125_ _07288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13312__I _07678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12909__A2 register_file\[18\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14426_ _01682_ register_file\[11\]\[9\] _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11638_ _06419_ _06623_ _06624_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13031__A1 _07455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14357_ _01611_ register_file\[6\]\[8\] _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11569_ _06579_ register_file\[11\]\[25\] _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11593__A1 _06375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16123__CLK clknet_leaf_288_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13308_ _07578_ _07634_ _07676_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14288_ _01800_ register_file\[1\]\[7\] _01801_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15323__A3 _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09538__A1 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16027_ _00415_ clknet_leaf_252_clk register_file\[6\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13334__A2 _07690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13239_ _07509_ _07632_ _07636_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16273__CLK clknet_leaf_158_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15087__A2 register_file\[22\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ _03134_ _03135_ _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08780_ _04095_ _04103_ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13098__A1 _07543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14834__A2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12845__A1 _07381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09710__A1 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09401_ _04576_ register_file\[19\]\[12\] _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14598__A1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09332_ _04644_ _04647_ _03796_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13270__A1 _07653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ _03799_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_178_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11820__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15011__A2 _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08214_ _03542_ _03543_ _03231_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08029__A1 _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13022__A1 _07491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09194_ _04508_ _04511_ _04094_ _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08145_ _03474_ _03150_ _03475_ _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08076_ _01111_ register_file\[25\]\[27\] _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11677__I _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13325__A2 register_file\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10139__A2 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11336__A1 _06440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08201__A1 _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11887__A2 register_file\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13892__I _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08978_ _03933_ register_file\[4\]\[6\] _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14825__A2 _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15640__CLK clknet_leaf_197_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13628__A3 _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12836__A1 _07381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07929_ _02929_ register_file\[9\]\[25\] _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09701__A1 _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10940_ _06189_ register_file\[2\]\[13\] _06190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10871_ _06131_ register_file\[30\]\[25\] _06141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15790__CLK clknet_leaf_127_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12610_ _07232_ _07233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13261__A1 _07646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12064__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13590_ _01110_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10075__A1 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12541_ _07190_ register_file\[22\]\[4\] _07192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15002__A2 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16146__CLK clknet_leaf_156_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13013__A1 _07484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15260_ _01104_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12472_ _07150_ register_file\[23\]\[8\] _07151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14211_ _01723_ _01724_ _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11423_ _06216_ _04219_ _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09766__B _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15191_ _02524_ register_file\[12\]\[18\] _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11575__A1 _06543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14142_ _01655_ _01656_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11354_ _06449_ _06454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11587__I _06593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16296__CLK clknet_leaf_80_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10305_ _03904_ _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_125_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13316__A2 register_file\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11285_ _06403_ register_file\[19\]\[14\] _06406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14073_ _01581_ _01588_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11327__A1 _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13024_ _07465_ _07494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_140_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10236_ _05338_ register_file\[13\]\[24\] _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11878__A2 _06778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09940__A1 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08896__I _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10167_ _05467_ _05470_ _05268_ _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10550__A2 register_file\[16\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12827__A1 _07257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14975_ _02230_ register_file\[27\]\[16\] _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10098_ _05399_ _05402_ _04183_ _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14292__A3 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12211__I _06068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13926_ _01443_ _01355_ _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10302__A2 register_file\[13\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13857_ _01351_ _01375_ _01195_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15241__A2 register_file\[24\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08259__A1 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12808_ _07362_ register_file\[1\]\[2\] _07365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13252__A1 _07522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12055__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16576_ _00964_ clknet_leaf_5_clk register_file\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13788_ _00998_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15527_ _01774_ _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12739_ _07318_ register_file\[20\]\[6\] _07324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11802__A2 register_file\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13042__I _07504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13004__A1 _07274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15458_ _00999_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13977__I _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14409_ _01916_ _01920_ _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12881__I _07407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15389_ _01055_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11566__A1 _06579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_292_clk clknet_5_5__leaf_clk clknet_leaf_292_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09950_ _05190_ register_file\[18\]\[20\] _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_3_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15663__CLK clknet_leaf_146_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08901_ _03923_ register_file\[1\]\[4\] _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09881_ _05187_ _05188_ _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_5_12__f_clk clknet_3_3_0_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11869__A2 register_file\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09931__A1 _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08832_ _03923_ register_file\[1\]\[3\] _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14807__A2 register_file\[26\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12818__A1 _07246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08763_ _03767_ register_file\[13\]\[3\] _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15480__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08498__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08694_ _04013_ _04016_ _04018_ _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15232__A2 register_file\[21\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16169__CLK clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12046__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13243__A1 _07638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09315_ _04499_ register_file\[3\]\[10\] _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09998__A1 _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14048__I _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09246_ _04560_ _04563_ _04078_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15588__B _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08670__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13887__I _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14743__A1 _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09177_ _04493_ _04495_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13546__A2 _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11557__A1 _06572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08128_ _03459_ register_file\[1\]\[27\] _01198_ _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_181_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08422__A1 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10525__B _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_283_clk clknet_5_5__leaf_clk clknet_leaf_283_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_107_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08973__A2 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08059_ _03222_ register_file\[17\]\[27\] _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11309__A1 _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput46 net46 rD[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__10780__A2 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput57 net57 rD[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11070_ _06268_ _06269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_103_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput68 net68 rD[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_163_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput79 net79 rS[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__12740__B _07324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10021_ _05323_ _05326_ _04452_ _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07834__B _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09605__I _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output58_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12809__A1 _07239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14274__A3 _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12031__I _06865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14760_ _02096_ register_file\[9\]\[13\] _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12285__A2 register_file\[31\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11972_ _06837_ register_file\[5\]\[13\] _06838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13482__A1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09150__A2 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13711_ _01081_ register_file\[28\]\[1\] _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10296__A1 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10923_ _06174_ register_file\[2\]\[6\] _06180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14691_ _02190_ _02199_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16430_ _00818_ clknet_leaf_147_clk register_file\[17\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13642_ register_file\[4\]\[0\] _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10854_ _06109_ register_file\[30\]\[22\] _06127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12037__A2 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09989__A1 _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16361_ _00749_ clknet_leaf_96_clk register_file\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14982__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13573_ _01093_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10785_ _06069_ _06052_ _06070_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11796__A1 _06658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10599__A2 _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15312_ _02812_ register_file\[26\]\[20\] _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12524_ _07034_ _07138_ _07180_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16292_ _00680_ clknet_leaf_74_clk register_file\[21\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08661__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15243_ _02743_ _02744_ _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12455_ _06965_ _07136_ _07140_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11548__A1 _06410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07795__I register_file\[3\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15686__CLK clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11406_ _06483_ register_file\[26\]\[24\] _06485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15174_ _02593_ register_file\[31\]\[18\] _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08413__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12386_ _06974_ _07098_ _07099_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10220__A1 _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14125_ _01639_ _01468_ _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_274_clk clknet_5_7__leaf_clk clknet_leaf_274_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11337_ _06159_ _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14056_ _01055_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11268_ _06391_ register_file\[19\]\[9\] _06394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13007_ _07454_ _07484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09913__A1 _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10219_ _05252_ register_file\[21\]\[24\] _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11199_ _06318_ _06348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10523__A2 register_file\[31\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14958_ register_file\[3\]\[15\] _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12276__A2 register_file\[31\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16311__CLK clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13909_ _01426_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14889_ _02394_ _02228_ _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12028__A2 _06864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13225__A1 _07583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16559_ _00947_ clknet_leaf_150_clk register_file\[29\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16461__CLK clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11787__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09100_ _04348_ register_file\[7\]\[7\] _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09031_ _04342_ _04351_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13528__A2 register_file\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13500__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12200__A2 _06976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_265_clk clknet_5_18__leaf_clk clknet_leaf_265_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_190_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08955__A2 register_file\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15150__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09933_ _05240_ _04973_ _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08707__A2 register_file\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09864_ _03831_ _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11711__A1 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09380__A2 register_file\[17\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08815_ _04077_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09795_ _04967_ register_file\[2\]\[17\] _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08746_ _03898_ register_file\[29\]\[2\] _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12267__A2 register_file\[31\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13464__A1 _07574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10278__A1 _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08677_ _03997_ _04000_ _04002_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08891__A1 _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14964__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10570_ _05864_ _05867_ _04873_ _05868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14716__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09229_ _04413_ register_file\[17\]\[9\] _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12240_ _07004_ _07000_ _07005_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08504__I _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_256_clk clknet_5_16__leaf_clk clknet_leaf_256_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12026__I _06865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12171_ _06911_ register_file\[3\]\[30\] _06956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11950__A1 _06652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11122_ _06297_ register_file\[27\]\[20\] _06301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11053_ _06139_ _06257_ _06258_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15930_ _00318_ clknet_leaf_256_clk register_file\[10\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14241__I _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16334__CLK clknet_leaf_145_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10004_ _05302_ _05310_ _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09371__A2 register_file\[8\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15861_ _00249_ clknet_leaf_218_clk register_file\[12\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14812_ _01986_ register_file\[29\]\[14\] _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14247__A3 _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15444__A2 register_file\[14\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15792_ _00180_ clknet_leaf_169_clk register_file\[19\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13455__A1 _07565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09123__A2 register_file\[30\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10269__A1 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14743_ _02164_ register_file\[19\]\[13\] _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11955_ _06822_ register_file\[5\]\[6\] _06828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15072__I _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10906_ _06166_ _06169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13207__A1 _07612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14674_ _02096_ register_file\[9\]\[12\] _02183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11886_ _06667_ _06785_ _06786_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16413_ _00801_ clknet_leaf_28_clk register_file\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13625_ _01021_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10837_ _06112_ _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16344_ _00732_ clknet_leaf_195_clk register_file\[20\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13556_ _01070_ _01073_ _01076_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12430__A2 register_file\[24\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10768_ _06042_ register_file\[30\]\[6\] _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14707__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12507_ _07134_ _07171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10441__A1 _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10944__I _06177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16275_ _00663_ clknet_leaf_209_clk register_file\[22\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13487_ net9 _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10699_ _05993_ _05994_ _05995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10992__A2 _06219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15226_ _02646_ register_file\[19\]\[19\] _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15380__A1 _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12438_ _07028_ _07126_ _07129_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12194__A1 _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_247_clk clknet_5_17__leaf_clk clknet_leaf_247_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15157_ _02650_ _02659_ _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12369_ _07087_ _07088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11941__A1 _06638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14108_ _01278_ register_file\[2\]\[5\] _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_138_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15132__A1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15088_ _01093_ _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14039_ _01554_ _01468_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12497__A2 _07160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I addrD[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09362__A2 _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15701__CLK clknet_leaf_211_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08600_ _03926_ _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_23_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09580_ _04892_ register_file\[21\]\[14\] _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13446__A1 _07555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08531_ _03839_ _03857_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15199__A1 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08462_ net5 _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08873__A1 _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15851__CLK clknet_leaf_122_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13749__A2 _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08393_ _03700_ _03720_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11015__I _06228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12421__A2 register_file\[24\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10432__A1 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09014_ _04312_ _04334_ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10983__A2 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12185__A1 _06965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_238_clk clknet_5_20__leaf_clk clknet_leaf_238_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08928__A2 register_file\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09050__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13921__A2 _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11932__A1 _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16357__CLK clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11685__I _06642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09916_ _05025_ register_file\[23\]\[19\] _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_8_clk_I clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10499__A1 _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09847_ _05090_ register_file\[16\]\[18\] _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09778_ _03765_ _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13437__A1 _07749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09105__A2 register_file\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08729_ _03870_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11999__A1 _06701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11740_ _06121_ _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14937__A1 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10671__A1 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11671_ _06032_ _06645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13410_ _07518_ _07738_ _07739_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_169_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10622_ _05668_ register_file\[31\]\[30\] _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14390_ _01564_ register_file\[29\]\[9\] _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12412__A2 _07112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13341_ _07694_ register_file\[29\]\[10\] _07698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10553_ _03871_ register_file\[19\]\[29\] _05851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10974__A2 _06206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16060_ _00448_ clknet_leaf_293_clk register_file\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13272_ _07641_ _07656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14165__A2 _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10484_ _03828_ register_file\[18\]\[28\] _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14680__B _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15011_ _02515_ _02270_ _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_229_clk clknet_5_21__leaf_clk clknet_leaf_229_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12223_ _06992_ _06988_ _06993_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09041__A1 _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11923__A1 _06803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15114__A1 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12154_ _06696_ _06943_ _06946_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11105_ _06290_ register_file\[27\]\[13\] _06291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15724__CLK clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12479__A2 register_file\[23\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12085_ _06899_ net30 _06905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13676__A1 _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09065__I _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11036_ _06108_ _06243_ _06248_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15913_ _00301_ clknet_leaf_111_clk register_file\[10\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15844_ _00232_ clknet_leaf_61_clk register_file\[12\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13428__A1 _07749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15874__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10939__I _06169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15775_ _00163_ clknet_leaf_12_clk register_file\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12987_ _07257_ _07466_ _07472_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12100__A1 _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13315__I _07681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14726_ _02229_ _02233_ _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11938_ _06814_ _06817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_45_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08855__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12651__A2 register_file\[21\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14657_ _01835_ register_file\[18\]\[12\] _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11869_ _06774_ register_file\[6\]\[4\] _06776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13608_ _01017_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08607__A1 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14588_ _02095_ _02097_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13600__A1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16327_ _00715_ clknet_leaf_80_clk register_file\[20\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10414__A1 _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13539_ _01059_ register_file\[25\]\[0\] _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09280__A1 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10965__A2 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16258_ _00646_ clknet_leaf_71_clk register_file\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15353__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07830__A2 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12167__A1 _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15209_ _02711_ _02378_ _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09032__A1 _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13903__A2 register_file\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16189_ _00577_ clknet_leaf_34_clk register_file\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11914__A1 _06696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10717__A2 register_file\[3\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11390__A2 _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14459__A3 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07962_ register_file\[3\]\[25\] _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_190_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09701_ _04992_ _05011_ _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07893_ _03226_ _01066_ _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11142__A2 register_file\[27\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15408__A2 register_file\[24\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09632_ _04926_ _04943_ _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13419__A1 _07529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09563_ _04859_ _04875_ _04876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09099__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08514_ _03840_ _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_70_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09494_ _04800_ _04807_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12642__A2 _07248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10653__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14919__A1 _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08445_ _03771_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15440__I _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14395__A2 register_file\[31\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08376_ _03703_ _03420_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14056__I _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08074__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15344__A1 _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07821__A2 register_file\[23\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12158__A1 _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15747__CLK clknet_leaf_54_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09023__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11905__A1 _06686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10708__A2 _06003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09574__A2 register_file\[18\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08377__A3 _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10533__B _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11381__A2 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12304__I _07049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15897__CLK clknet_leaf_261_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09326__A2 register_file\[25\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12330__A1 _06999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12910_ _07259_ _07425_ _07426_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13890_ _01402_ _01407_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_171_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12841_ _07381_ register_file\[1\]\[15\] _07385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10759__I _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10892__A1 _06156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_261_clk_I clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14083__A1 _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15560_ _02889_ register_file\[24\]\[23\] _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12772_ _07321_ _07343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__A1 _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14511_ _01688_ register_file\[12\]\[10\] _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11723_ _06099_ _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10644__A1 _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15491_ _02986_ _02989_ _02658_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14442_ _01530_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_276_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11654_ _06436_ _06630_ _06633_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12397__A1 _07102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10605_ _05900_ _05901_ _05902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14373_ _01800_ register_file\[1\]\[8\] _01801_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11585_ _06591_ _06592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10947__A2 register_file\[2\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16112_ _00500_ clknet_leaf_226_clk register_file\[3\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13324_ _07513_ _07680_ _07687_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15335__A1 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10536_ _05640_ register_file\[1\]\[28\] _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12149__A1 _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16043_ _00431_ clknet_leaf_289_clk register_file\[5\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13255_ _07633_ _07646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10467_ _05565_ register_file\[24\]\[27\] _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13897__A1 _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12206_ _06980_ _06976_ _06981_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09565__A2 register_file\[8\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13186_ _07536_ _07601_ _07604_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10398_ _05689_ _05698_ _05699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12214__I _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12137_ _06933_ register_file\[3\]\[15\] _06937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_214_clk_I clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09317__A2 register_file\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14310__A2 register_file\[31\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12068_ _06873_ _06895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_46_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12321__A1 _07054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11124__A2 register_file\[27\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11019_ _06078_ _06236_ _06238_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07879__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09523__I _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12872__A2 _07398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_229_clk_I clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15827_ _00215_ clknet_leaf_173_clk register_file\[26\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16052__CLK clknet_leaf_230_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15758_ _00146_ clknet_leaf_148_clk register_file\[13\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12624__A2 _07233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10635__A1 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14709_ _01370_ _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15689_ _00077_ clknet_leaf_101_clk register_file\[28\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15260__I _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08230_ _01090_ register_file\[26\]\[29\] _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15574__A1 _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12388__A1 _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08161_ _01135_ register_file\[21\]\[28\] _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10938__A2 _06185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11060__A1 _06218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15326__A1 _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08092_ _03415_ _03423_ _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09005__A1 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13888__A1 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08602__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10353__B _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12560__A1 _06990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12124__I _06921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08994_ _04313_ _04314_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14301__A2 register_file\[27\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07945_ _01051_ _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12312__A1 _07054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11115__A2 _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07876_ _03209_ _03210_ _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12863__A2 _07391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09433__I _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09615_ _04727_ register_file\[13\]\[15\] _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _04849_ _04858_ _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_5_28__f_clk_I clknet_3_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08819__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16545__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10626__A1 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09477_ _04789_ _04790_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15170__I _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07888__I _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08428_ _03755_ _01182_ _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14368__A2 register_file\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12379__A1 _07094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09244__A1 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08359_ _00995_ _03686_ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13040__A2 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10929__A2 _06178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11370_ _06462_ register_file\[26\]\[9\] _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09795__A2 register_file\[2\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10321_ _05425_ register_file\[24\]\[25\] _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14514__I _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09547__A2 register_file\[29\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13040_ _06216_ _03854_ _07503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output88_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10252_ _05423_ register_file\[25\]\[24\] _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10183_ _05418_ register_file\[7\]\[23\] _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14991_ _02495_ _02331_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11106__A2 _06286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13942_ _01458_ _01459_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12854__A2 _07391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11094__B _06284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10865__A1 _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13873_ _01043_ register_file\[22\]\[3\] _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_80_clk_I clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15612_ _00000_ clknet_leaf_37_clk register_file\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12824_ _07374_ register_file\[1\]\[8\] _07375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16592_ _00980_ clknet_leaf_176_clk register_file\[9\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12606__A2 _07186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15543_ register_file\[5\]\[22\] _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10617__A1 _05906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12755_ _07313_ _07333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09483__A1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15912__CLK clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11290__A1 _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11706_ _06077_ _06670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10093__A2 register_file\[28\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14359__A2 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15474_ _02927_ _02973_ _02888_ net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12686_ _07286_ _07284_ _07287_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_95_clk_I clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14425_ _01936_ _01855_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11637_ _06620_ register_file\[10\]\[20\] _06624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13031__A2 register_file\[17\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11042__A1 _06247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14356_ _01861_ _01868_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11568_ _06553_ _06582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12790__A1 _07300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13307_ _07631_ register_file\[14\]\[30\] _07676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11593__A2 _06592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10519_ _05756_ register_file\[29\]\[28\] _05818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14287_ _01370_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11499_ _06495_ register_file\[12\]\[30\] _06540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09518__I _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16026_ _00414_ clknet_leaf_252_clk register_file\[6\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09538__A2 register_file\[24\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13238_ _07634_ register_file\[14\]\[1\] _07636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_153_clk_I clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12542__A1 _06972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16418__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09962__B _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13169_ _07590_ register_file\[15\]\[5\] _07595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08210__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_33_clk_I clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14295__A1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13098__A2 _07544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_168_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12845__A2 register_file\[1\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_48_clk_I clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14047__A1 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09400_ _04441_ register_file\[18\]\[12\] _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14598__A2 register_file\[12\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09331_ _04645_ _04646_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08277__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09262_ _04574_ _04578_ _03943_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08213_ _03229_ register_file\[18\]\[29\] _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09226__A1 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09193_ _04509_ _04510_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12119__I _06913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08029__A2 register_file\[15\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13022__A2 register_file\[17\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11033__A1 _06104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08144_ _03235_ register_file\[29\]\[28\] _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07788__A1 _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12781__A1 _07290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10862__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08075_ _03243_ register_file\[24\]\[27\] _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11179__B _06336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16098__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12533__A1 _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11336__A2 _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ _04265_ _04297_ _04298_ net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07928_ _03181_ register_file\[8\]\[25\] _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12836__A2 register_file\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07859_ _02857_ register_file\[14\]\[24\] _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15935__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10870_ _06051_ _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_147_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14589__A2 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12738__B _07323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09529_ _04826_ _04842_ _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09465__A1 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13261__A2 register_file\[14\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10075__A2 register_file\[17\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11272__A1 _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12540_ _06969_ _07184_ _07191_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10258__B _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12471_ _07137_ _07150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09217__A1 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13013__A2 register_file\[17\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14210__A1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14210_ _01550_ register_file\[25\]\[7\] _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11024__A1 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11422_ _06444_ _06450_ _06493_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15190_ _02688_ _02692_ _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09768__A2 _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07779__A1 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10772__I _06059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14141_ _01308_ register_file\[17\]\[6\] _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14244__I _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11353_ _06375_ _06448_ _06453_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ _05604_ _05605_ _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14513__A2 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14072_ _01584_ _01587_ _01237_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11284_ _06090_ _06405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12524__A1 _07034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11327__A2 _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13023_ _07293_ _07487_ _07493_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10235_ _05534_ _05537_ _05268_ _05538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15069__A3 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09940__A2 register_file\[30\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10166_ _05468_ _05469_ _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12827__A2 _07370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14974_ _02478_ _02228_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10097_ _05400_ _05401_ _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10838__A1 _06109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13925_ register_file\[7\]\[3\] _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13856_ _01364_ _01374_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12807_ _07237_ _07360_ _07364_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09456__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13787_ _01056_ register_file\[24\]\[2\] _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08259__A2 register_file\[6\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16575_ _00963_ clknet_leaf_5_clk register_file\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13252__A2 _07642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10999_ _06041_ _06219_ _06226_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12738_ _07246_ _07322_ _07323_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15526_ _02940_ register_file\[12\]\[22\] _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15529__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09208__A1 _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15457_ register_file\[5\]\[21\] _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12669_ _07274_ _07272_ _07275_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13004__A2 _07480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08861__B _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14408_ _01917_ _01918_ _01919_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14752__A2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15388_ _02844_ _02887_ _02888_ net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11778__I _06718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12763__A1 _07333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11566__A2 register_file\[11\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16240__CLK clknet_leaf_151_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14339_ _01850_ _01851_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15808__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12515__A1 _07171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16009_ _00397_ clknet_leaf_292_clk register_file\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08900_ _04154_ register_file\[3\]\[4\] _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09880_ _04919_ register_file\[24\]\[19\] _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16390__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ _04154_ register_file\[3\]\[3\] _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09931__A2 register_file\[1\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14268__A1 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10631__B _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08762_ _04048_ _04086_ _03936_ net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12818__A2 _07370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08101__B _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08693_ _04017_ _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13491__A2 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13243__A2 register_file\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13233__I _07631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09314_ _04630_ register_file\[2\]\[10\] _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09998__A2 register_file\[3\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14991__A2 _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09245_ _04561_ _04562_ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08670__A2 register_file\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08771__B _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11006__A1 _06225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09176_ _04494_ register_file\[15\]\[8\] _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12754__A1 _07264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ _01005_ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_179_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08422__A2 register_file\[22\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08058_ _03306_ register_file\[16\]\[27\] _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12506__A1 _07016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11309__A2 register_file\[19\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput47 net47 rD[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput58 net58 rD[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_150_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput69 net69 rD[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08186__A1 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10020_ _05324_ _05325_ _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14259__A1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10541__B _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13408__I _07737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07933__A1 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12809__A2 _07360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11971_ _06817_ _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09686__A1 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13482__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13710_ _01226_ _01229_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10922_ _06050_ _06178_ _06179_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10296__A2 register_file\[8\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11493__A1 _06531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14690_ _02195_ _02198_ _02030_ _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16113__CLK clknet_leaf_226_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13641_ _01161_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10853_ _06125_ _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09438__A1 _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10767__I _06055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14431__A1 _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16360_ _00748_ clknet_leaf_82_clk register_file\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09989__A2 register_file\[21\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13572_ _01092_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10784_ _06065_ register_file\[30\]\[9\] _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14982__A2 register_file\[30\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13785__A3 _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15311_ _01042_ _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12993__A1 _07470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12523_ _07135_ register_file\[23\]\[30\] _07180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11796__A2 _06730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16291_ _00679_ clknet_leaf_68_clk register_file\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09777__B _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08661__A2 register_file\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15242_ _02576_ register_file\[25\]\[19\] _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12454_ _07138_ register_file\[23\]\[1\] _07140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12745__A1 _07254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11548__A2 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11405_ _06426_ _06479_ _06484_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15173_ _02590_ register_file\[30\]\[18\] _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12385_ _07094_ register_file\[24\]\[5\] _07099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09610__A1 _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08413__A2 register_file\[16\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14124_ _01638_ _01553_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10220__A2 register_file\[20\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11336_ _06440_ _06432_ _06441_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14055_ _01562_ _01570_ _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11267_ _06068_ _06393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13006_ _07276_ _07480_ _07483_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13170__A1 _07518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10218_ _05517_ _05520_ _04018_ _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09913__A2 register_file\[20\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11198_ _06104_ _06344_ _06347_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10149_ _05452_ register_file\[30\]\[23\] _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09677__A1 _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14957_ _02131_ register_file\[2\]\[15\] _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14670__A1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11484__A1 _06531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13908_ net9 _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14888_ _02392_ _02393_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09429__A1 _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13839_ register_file\[4\]\[2\] _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14422__A1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13225__A2 register_file\[15\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14973__A2 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16558_ _00946_ clknet_leaf_150_clk register_file\[29\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13988__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12984__A1 _07470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15509_ _03007_ register_file\[30\]\[22\] _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16489_ _00877_ clknet_leaf_110_clk register_file\[15\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09030_ _04345_ _04350_ _04068_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15630__CLK clknet_leaf_152_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11301__I _06112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14489__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09932_ _05237_ _05238_ _05239_ _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14612__I register_file\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07935__B _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15150__A2 register_file\[21\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13161__A1 _07511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09863_ _04967_ register_file\[2\]\[18\] _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07915__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11711__A2 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08814_ _04136_ _04137_ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _05100_ _05103_ _04220_ _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08745_ _04058_ _04069_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09668__A1 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14661__A1 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11971__I _06817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13464__A2 _07766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11475__A1 _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10278__A2 register_file\[16\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08676_ _04001_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_81_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09441__I _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14413__A1 _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11227__A1 _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13767__A3 _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09840__A1 _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09228_ _04542_ _04545_ _04118_ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14716__A2 register_file\[24\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12727__A1 _07237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09159_ _04476_ _04477_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11211__I _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12170_ _06712_ _06950_ _06955_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11121_ _06278_ _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11950__A2 _06816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14522__I _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15141__A2 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output70_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11052_ _06254_ register_file\[28\]\[25\] _06258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10003_ _05308_ _05309_ _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15860_ _00248_ clknet_leaf_175_clk register_file\[12\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14811_ _01035_ _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15791_ _00179_ clknet_leaf_127_clk register_file\[19\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09659__A1 _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13455__A2 _07759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11466__A1 _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10269__A2 register_file\[2\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14742_ _02248_ _02249_ _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11954_ _06654_ _06826_ _06827_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09351__I _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10905_ _06167_ _06168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14673_ _01932_ register_file\[8\]\[12\] _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13207__A2 register_file\[15\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_192_clk clknet_5_25__leaf_clk clknet_leaf_192_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11885_ _06782_ register_file\[6\]\[10\] _06786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13624_ _01140_ _01141_ _01144_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11218__A1 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16412_ _00800_ clknet_leaf_277_clk register_file\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10836_ _06111_ _06112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15653__CLK clknet_leaf_69_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14955__A2 _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12966__A1 _07458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15302__B _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16343_ _00731_ clknet_leaf_197_clk register_file\[20\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13555_ _01075_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10767_ _06055_ _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09831__A1 _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12506_ _07016_ _07167_ _07170_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16274_ _00662_ clknet_leaf_158_clk register_file\[22\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10441__A2 register_file\[14\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13486_ _01002_ _01006_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10698_ _05752_ register_file\[7\]\[31\] _05994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12718__A1 _07308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15225_ _02726_ _01292_ _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12437_ _07123_ register_file\[24\]\[27\] _07129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11121__I _06278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08398__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13391__A1 _06316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15156_ _02654_ _02657_ _02658_ _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_5_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12368_ _07086_ _07087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15528__I _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14107_ _01176_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11319_ _06427_ register_file\[19\]\[24\] _06430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11941__A2 _06816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15087_ _02590_ register_file\[22\]\[17\] _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15132__A2 register_file\[1\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12299_ _07046_ register_file\[25\]\[3\] _07047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16159__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13143__A1 _07504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14038_ _01552_ _01553_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13694__A2 _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13446__A2 _07759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15989_ _00377_ clknet_leaf_233_clk register_file\[7\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11791__I _06721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08530_ _03846_ _03853_ _03856_ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11457__A1 _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ _03781_ _03787_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15199__A2 register_file\[6\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_183_clk clknet_5_28__leaf_clk clknet_leaf_183_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08873__A2 register_file\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11209__A1 _06348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08392_ _03712_ _03719_ _01505_ _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12957__A1 _07407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09822__A1 _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10432__A2 register_file\[8\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09013_ _04324_ _04333_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12709__A1 _07302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08389__A1 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12185__A2 _06961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13382__A1 _07572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10870__I _06051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11932__A2 _06770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14342__I _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13134__A1 _07563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09915_ _05023_ register_file\[22\]\[19\] _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09889__A1 _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14882__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09846_ _05088_ register_file\[17\]\[18\] _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10499__A2 register_file\[6\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08561__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09777_ _05081_ _05086_ _04057_ _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11448__A1 _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08728_ _04052_ register_file\[6\]\[2\] _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15676__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11999__A2 _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08659_ _03983_ _03984_ _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_174_clk clknet_5_29__leaf_clk clknet_leaf_174_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_14_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11670_ _06638_ _06641_ _06644_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14937__A2 register_file\[14\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12948__A1 _07298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10621_ _05666_ register_file\[30\]\[30\] _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09813__A1 _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13340_ _07689_ _07697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11620__A1 _06613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10552_ _03868_ register_file\[18\]\[29\] _05850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14961__B _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13271_ _07541_ _07649_ _07655_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10483_ _05780_ _05781_ _05782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15010_ _02512_ _02514_ _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12222_ _06983_ register_file\[31\]\[12\] _06993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13373__A1 _07562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12176__A2 _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__A1 _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09041__A2 register_file\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11923__A2 register_file\[6\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12153_ _06940_ register_file\[3\]\[22\] _06946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13125__A1 _07562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11104_ _06270_ _06290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12084_ _03371_ _06902_ _06904_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14873__A1 _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13676__A2 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11035_ _06247_ register_file\[28\]\[18\] _06248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15912_ _00300_ clknet_leaf_109_clk register_file\[10\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16451__CLK clknet_leaf_56_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11687__A1 _06650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15843_ _00231_ clknet_leaf_56_clk register_file\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14625__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12500__I _07145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12986_ _07470_ register_file\[17\]\[9\] _07472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15774_ _00162_ clknet_leaf_29_clk register_file\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12100__A2 register_file\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14725_ _02231_ _02232_ _01982_ _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_165_clk clknet_5_31__leaf_clk clknet_leaf_165_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11937_ _06815_ _06816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11116__I _06267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08855__A2 register_file\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14656_ _02164_ register_file\[19\]\[12\] _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14928__A2 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11868_ _06649_ _06768_ _06775_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10819_ net18 _06098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13607_ _01118_ _01127_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_186_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09804__A1 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14587_ _02096_ register_file\[9\]\[11\] _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11799_ _06721_ _06734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08607__A2 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16326_ _00714_ clknet_leaf_81_clk register_file\[20\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11611__A1 _06393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09030__B _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13538_ _01058_ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09280__A2 register_file\[17\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16257_ _00645_ clknet_leaf_71_clk register_file\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13469_ _07727_ register_file\[9\]\[31\] _07773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12167__A2 register_file\[3\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15208_ _02705_ _02710_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09032__A2 register_file\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16188_ _00576_ clknet_leaf_35_clk register_file\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10178__A1 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11786__I _06721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11914__A2 _06799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15139_ _02390_ register_file\[17\]\[18\] _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08791__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ _02964_ register_file\[2\]\[25\] _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09700_ _05001_ _05010_ _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07892_ _03224_ _03225_ _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09631_ _04933_ _04942_ _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13419__A2 _07738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10350__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09562_ _04866_ _04874_ _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09099__A2 register_file\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08513_ _03798_ _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_24_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09493_ _04803_ _04806_ _04400_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10102__A1 _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_156_clk clknet_5_30__leaf_clk clknet_leaf_156_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08444_ _03770_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__14919__A2 register_file\[23\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11850__A1 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08375_ register_file\[9\]\[31\] _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11602__A1 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16324__CLK clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15344__A2 register_file\[8\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13355__A1 _07701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10169__A1 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09023__A2 register_file\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11696__I _06642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11905__A2 _06792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16474__CLK clknet_leaf_253_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13107__A1 _07551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08782__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14855__A1 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11669__A1 _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12330__A2 _07064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09829_ _05004_ register_file\[8\]\[18\] _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14607__A1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12840_ _07369_ _07384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10892__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15280__A1 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12771_ _07281_ _07336_ _07342_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_147_clk clknet_5_27__leaf_clk clknet_leaf_147_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13830__A2 _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14510_ _02017_ _02020_ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11722_ _06679_ _06680_ _06681_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15490_ _02987_ _02738_ _02988_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10644__A2 register_file\[22\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11841__A1 _06755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14441_ _01950_ _01952_ _01702_ _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10775__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11653_ _06627_ register_file\[10\]\[27\] _06633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15583__A2 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12397__A2 register_file\[24\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10604_ _03824_ register_file\[8\]\[30\] _05901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14372_ _01623_ _01881_ _01884_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11584_ _06590_ _06591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16111_ _00499_ clknet_leaf_190_clk register_file\[3\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13323_ _07686_ register_file\[29\]\[3\] _07687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _03832_ register_file\[3\]\[28\] _05834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15335__A2 register_file\[20\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14138__A3 _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13346__A1 _07536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12149__A2 register_file\[3\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13254_ _07524_ _07642_ _07645_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16042_ _00430_ clknet_leaf_289_clk register_file\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10466_ _05563_ register_file\[25\]\[27\] _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09014__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13897__A2 register_file\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12205_ _06970_ register_file\[31\]\[7\] _06981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13185_ _07598_ register_file\[15\]\[12\] _07604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10397_ _05692_ _05697_ _03992_ _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08773__A1 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12136_ _06921_ _06936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15841__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10580__A1 _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12067_ _02787_ _06888_ _06894_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08525__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12321__A2 register_file\[25\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ _06233_ register_file\[28\]\[11\] _06238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10332__A1 _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15826_ _00214_ clknet_leaf_169_clk register_file\[26\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_138_clk clknet_5_26__leaf_clk clknet_leaf_138_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15757_ _00145_ clknet_leaf_148_clk register_file\[13\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12969_ _07239_ _07456_ _07461_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14708_ _01185_ _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11832__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15688_ _00076_ clknet_leaf_84_clk register_file\[28\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15023__A1 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14639_ _02146_ _02147_ _01982_ _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15574__A2 register_file\[30\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14377__A3 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13061__I _07506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12388__A2 _07098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08160_ _01130_ register_file\[20\]\[28\] _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08056__A3 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_7_clk_I clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10399__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16309_ _00697_ clknet_leaf_206_clk register_file\[21\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15326__A2 register_file\[16\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16497__CLK clknet_leaf_175_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08091_ _03418_ _03422_ _03340_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11060__A2 register_file\[28\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_310_clk clknet_5_1__leaf_clk clknet_leaf_310_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_173_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07803__A3 _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13337__A1 _07526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09005__A2 register_file\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13888__A2 register_file\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11899__A1 _06789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08764__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12560__A2 _07201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08993_ _04031_ register_file\[16\]\[6\] _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07944_ _03275_ _02945_ _03277_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09714__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12312__A2 register_file\[25\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07875_ _01021_ _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10323__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09614_ _04916_ _04925_ _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09545_ _04852_ _04857_ _04382_ _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_129_clk clknet_5_27__leaf_clk clknet_leaf_129_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15451__I register_file\[7\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09476_ _04518_ register_file\[27\]\[13\] _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10626__A2 register_file\[16\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15014__A1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08295__A3 _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08427_ register_file\[21\]\[31\] _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15714__CLK clknet_leaf_54_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12379__A2 register_file\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08358_ register_file\[4\]\[31\] _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09244__A2 register_file\[31\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08289_ _01081_ register_file\[20\]\[30\] _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_301_clk clknet_5_4__leaf_clk clknet_leaf_301_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10320_ _05423_ register_file\[25\]\[25\] _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15864__CLK clknet_leaf_260_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10251_ _05550_ _05553_ _05421_ _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08755__A1 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10182_ _05416_ register_file\[6\]\[23\] _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14828__A1 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14990_ _02493_ _02494_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13941_ _01369_ register_file\[1\]\[3\] _01371_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10314__A1 _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10865__A2 register_file\[30\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13872_ _01388_ _01036_ _01389_ _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15253__A1 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15611_ _03106_ _03107_ _03108_ _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12823_ _07361_ _07374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16591_ _00979_ clknet_leaf_189_clk register_file\[9\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15361__I _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13803__A2 _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15542_ _02786_ _03040_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11814__A1 _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12754_ _07264_ _07329_ _07332_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09483__A2 register_file\[18\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11705_ _06667_ _06668_ _06669_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12685_ _07279_ register_file\[21\]\[21\] _07287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11290__A2 _06408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15473_ _02949_ _02972_ _02886_ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14424_ _01935_ _01853_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11636_ _06601_ _06623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_50_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11042__A2 register_file\[28\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15308__A2 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14355_ _01864_ _01867_ _01608_ _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14705__I register_file\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11567_ _06429_ _06575_ _06581_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_183_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13319__A1 _07509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07797__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12790__A2 _07350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13306_ _07576_ _07670_ _07675_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10518_ _05813_ _05816_ _04118_ _05817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14286_ _01185_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11498_ _06440_ _06534_ _06539_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16025_ _00413_ clknet_leaf_243_clk register_file\[6\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13237_ _07502_ _07632_ _07635_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12225__I _06962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10449_ _05747_ _05748_ _05749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14531__A3 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08746__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12542__A2 _07184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13168_ _07593_ _07594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10553__A1 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12119_ _06913_ _06926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13099_ _06098_ _07546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14295__A2 register_file\[25\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__A1 _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14047__A2 register_file\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15809_ _00197_ clknet_leaf_50_clk register_file\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12895__I _07409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09330_ _04576_ register_file\[27\]\[11\] _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11805__A1 _06734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _04575_ _04577_ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15547__A2 _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11304__I _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08212_ _01069_ register_file\[19\]\[29\] _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09192_ _04233_ register_file\[15\]\[9\] _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15887__CLK clknet_leaf_186_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08143_ _01081_ register_file\[28\]\[28\] _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12230__A1 _06997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11033__A2 _06243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15220__B _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14615__I _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08985__A1 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12781__A2 _07343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08074_ _03398_ _03405_ _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_260_clk_I clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08737__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12533__A2 _07184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13730__A1 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08976_ _03935_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_25_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input32_I new_value[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_275_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16512__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12297__A1 _06967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07927_ _03242_ _03260_ _03179_ _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_151_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09162__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07858_ _03191_ _03026_ _03192_ _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15235__A1 _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14038__A2 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12049__A1 _06878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07789_ register_file\[5\]\[23\] _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09528_ _04835_ _04841_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09459_ _04771_ _04772_ _04773_ _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_213_clk_I clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13549__A1 _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12470_ _06980_ _07146_ _07149_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11421_ _06447_ register_file\[26\]\[31\] _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11024__A2 _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07779__A2 register_file\[15\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14140_ _01572_ register_file\[16\]\[6\] _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11352_ _06450_ register_file\[26\]\[2\] _06453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_228_clk_I clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16042__CLK clknet_leaf_289_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10303_ _05340_ register_file\[12\]\[25\] _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14071_ _01585_ _01326_ _01586_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_153_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11283_ _06402_ _06396_ _06404_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13022_ _07491_ register_file\[17\]\[24\] _07493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08728__A1 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12524__A2 _07138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13721__A1 _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10234_ _05535_ _05536_ _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10535__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11884__I _06777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15356__I _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10165_ _05334_ register_file\[11\]\[23\] _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16192__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15474__A1 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07951__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14973_ _02477_ _02393_ _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10096_ _05334_ register_file\[31\]\[22\] _05401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09153__A1 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13924_ _01152_ register_file\[6\]\[3\] _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_43_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15226__A1 _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08900__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13855_ _01373_ _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13604__I _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12806_ _07362_ register_file\[1\]\[1\] _07364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16574_ _00962_ clknet_leaf_305_clk register_file\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09456__A2 register_file\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13786_ _01297_ _01304_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10998_ _06225_ register_file\[28\]\[3\] _06226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15525_ _03020_ _03023_ _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12737_ _07318_ register_file\[20\]\[5\] _07323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15529__A2 register_file\[13\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12460__A1 _06969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15456_ _02786_ _02955_ _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12668_ _07267_ register_file\[21\]\[16\] _07275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14201__A2 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14407_ _01075_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10963__I _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12212__A1 _06983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11619_ _06593_ _06613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15387_ _01199_ _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12599_ _07183_ register_file\[22\]\[28\] _07226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08967__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12763__A2 register_file\[20\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14338_ _01676_ register_file\[9\]\[8\] _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10774__A1 _06060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08431__A3 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14269_ _01772_ _01782_ _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12515__A2 register_file\[23\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13712__A1 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16008_ _00396_ clknet_leaf_296_clk register_file\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16535__CLK clknet_leaf_226_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09392__A1 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ _03919_ _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15465__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12279__A1 _06960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08761_ _04070_ _04085_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09144__A1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08692_ _03854_ _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15215__B _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13514__I _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13779__A1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08608__I _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ _03916_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14440__A2 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11034__I _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_60_clk clknet_5_8__leaf_clk clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09244_ _04494_ register_file\[31\]\[9\] _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16065__CLK clknet_leaf_313_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12203__A1 _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09175_ _04148_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11006__A2 register_file\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10873__I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09439__I _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08126_ _03294_ _03455_ _03457_ _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12754__A2 _07329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08057_ _03343_ _03389_ _03305_ net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12506__A2 _07167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput48 net48 rD[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_143_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput59 net59 rD[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_118_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09383__A1 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08186__A2 register_file\[6\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15902__CLK clknet_leaf_303_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11190__A1 _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15456__A1 _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07933__A2 register_file\[11\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_94_clk_I clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08959_ _04211_ register_file\[5\]\[5\] _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10113__I _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11970_ _06672_ _06833_ _06836_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10921_ _06174_ register_file\[2\]\[5\] _06179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11493__A2 register_file\[12\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13640_ _00993_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10852_ _06124_ _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_5_12__f_clk_I clknet_3_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14431__A2 register_file\[13\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_152_clk_I clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10783_ _06068_ _06069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12442__A1 _07032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13571_ _01023_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16408__CLK clknet_leaf_195_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15310_ _02646_ register_file\[27\]\[20\] _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12993__A2 register_file\[17\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12522_ _07032_ _07174_ _07179_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_32_clk_I clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16290_ _00678_ clknet_leaf_68_clk register_file\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11879__I _06769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10783__I _06068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15241_ _02411_ register_file\[24\]\[19\] _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12453_ _06958_ _07136_ _07139_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_167_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12745__A2 _07322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11404_ _06483_ register_file\[26\]\[23\] _06484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12384_ _07097_ _07098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15172_ _02671_ _02672_ _02674_ _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__16558__CLK clknet_leaf_150_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09610__A2 register_file\[18\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10756__A1 _06042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_47_clk_I clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14123_ _01636_ _01637_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11335_ _06368_ register_file\[19\]\[29\] _06441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14498__A2 _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11266_ _06390_ _06384_ _06392_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14054_ _01566_ _01569_ _01395_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15086__I _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__A1 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13005_ _07477_ register_file\[17\]\[17\] _07483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10217_ _05518_ _05519_ _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13170__A2 _07594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11197_ _06341_ register_file\[13\]\[17\] _06347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11181__A1 _06334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__A2 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10148_ _03827_ _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_105_clk_I clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10079_ _05248_ register_file\[19\]\[22\] _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14956_ _01176_ _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09677__A2 register_file\[22\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13907_ _01422_ _01424_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14887_ _01062_ _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13838_ _01352_ _01356_ _01266_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14422__A2 register_file\[9\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16557_ _00945_ clknet_leaf_129_clk register_file\[29\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12433__A1 _07123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13769_ _01202_ register_file\[16\]\[2\] _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_42_clk clknet_5_12__leaf_clk clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_189_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15508_ _01122_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12984__A2 register_file\[17\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16488_ _00876_ clknet_leaf_48_clk register_file\[15\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10995__A1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07860__A1 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15439_ _02933_ _02938_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09259__I _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09931_ _04970_ register_file\[1\]\[19\] _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13161__A2 _07584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ _05165_ _05170_ _04068_ _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11172__A1 _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08813_ _03988_ register_file\[31\]\[3\] _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _05101_ _05102_ _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08744_ _04063_ _04066_ _04068_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09668__A2 register_file\[24\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14661__A2 register_file\[20\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10868__I _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08675_ _03893_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12672__A1 _07276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11475__A2 _06520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__A2 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14413__A2 register_file\[22\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12424__A1 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09878__B _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_33_clk clknet_5_6__leaf_clk clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_50_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11699__I _06068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10986__A1 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14177__A1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09227_ _04543_ _04544_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09158_ _04409_ register_file\[11\]\[8\] _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13924__A1 _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12727__A2 _07312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08109_ _03439_ _03361_ _03440_ _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09089_ _03870_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11120_ _06113_ _06293_ _06299_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08801__I _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09356__A1 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11051_ _06228_ _06257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_1_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12323__I _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09118__B _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output63_I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11163__A1 _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10002_ _04636_ _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07906__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10910__A1 _06170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08957__B _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09108__A1 _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14810_ _02235_ register_file\[28\]\[14\] _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14101__A1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15790_ _00178_ clknet_leaf_127_clk register_file\[19\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09659__A2 register_file\[1\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10778__I _06028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14741_ _01008_ _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11466__A2 _06520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11953_ _06822_ register_file\[5\]\[5\] _06827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16230__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13154__I _07582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10904_ _06166_ _06167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14672_ _02157_ _02180_ _01930_ _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11884_ _06777_ _06785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_45_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14404__A2 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15601__A1 _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16411_ _00799_ clknet_leaf_277_clk register_file\[18\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13623_ _01143_ register_file\[15\]\[0\] _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10835_ net21 _06111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11218__A2 _06358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_24_clk clknet_5_3__leaf_clk clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16342_ _00730_ clknet_leaf_182_clk register_file\[20\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08095__A1 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13554_ _01074_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10766_ _06054_ _06055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16380__CLK clknet_leaf_278_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09831__A2 register_file\[10\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10977__A1 _06167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14168__A1 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12505_ _07164_ register_file\[23\]\[22\] _07170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16273_ _00661_ clknet_leaf_158_clk register_file\[22\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15948__CLK clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10697_ _05750_ register_file\[6\]\[31\] _05993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13485_ _01005_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_173_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15224_ _02725_ _02393_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12718__A2 _07235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12436_ _07026_ _07126_ _07128_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15155_ _01100_ _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13391__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12367_ _04067_ _06215_ _07086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14106_ _01621_ _01538_ _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11318_ _06134_ _06429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15086_ _01089_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12298_ _07041_ _07046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13143__A2 register_file\[16\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14037_ _01005_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11249_ _06045_ _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10901__A1 _06026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15988_ _00376_ clknet_leaf_229_clk register_file\[7\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09542__I _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14643__A2 _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12654__A1 _07255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14939_ _02444_ register_file\[15\]\[15\] _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08460_ _03786_ register_file\[27\]\[0\] _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12406__A1 _07109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11209__A2 register_file\[13\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08391_ _03715_ _03718_ _01173_ _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_15_clk clknet_5_2__leaf_clk clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08086__A1 _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12957__A2 register_file\[18\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12408__I _07097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09012_ _04329_ _04332_ _04262_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12709__A2 _07296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08389__A2 register_file\[15\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13382__A2 _07718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14623__I register_file\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11393__A1 _06414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15123__A3 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14331__A1 _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09914_ _05220_ _05221_ _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12143__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13134__A2 register_file\[16\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11145__A1 _06160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09889__A2 register_file\[5\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09845_ _05150_ _05153_ _04675_ _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12893__A1 _07414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16253__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _05083_ _05085_ _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08727_ _03867_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12645__A1 _07257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11448__A2 register_file\[12\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08658_ _03883_ register_file\[20\]\[1\] _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output101_I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08589_ _03806_ _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_42_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10620_ _05915_ _05916_ _05917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12948__A2 _07446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13070__A1 _07524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10959__A1 _06196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09813__A2 register_file\[5\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07824__A1 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10551_ _05847_ _05848_ _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11620__A2 register_file\[10\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13270_ _07653_ register_file\[14\]\[14\] _07655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13858__B _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10482_ _03824_ register_file\[16\]\[28\] _05781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15362__A3 _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12221_ _06081_ _06992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13373__A2 _07711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09627__I _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12152_ _06694_ _06943_ _06945_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11103_ _06082_ _06286_ _06289_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09329__A1 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13125__A2 _07556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12083_ _06899_ net29 _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11136__A1 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15911_ _00299_ clknet_leaf_109_clk register_file\[10\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14873__A2 register_file\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11034_ _06217_ _06247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08001__A1 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12988__I _07465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11687__A2 register_file\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12884__A1 _07410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15364__I _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15842_ _00230_ clknet_leaf_52_clk register_file\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15620__CLK clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15773_ _00161_ clknet_leaf_280_clk register_file\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12985_ _07254_ _07466_ _07471_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09501__A1 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14724_ _01980_ register_file\[26\]\[13\] _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11936_ _06814_ _06815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_166_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14655_ _01119_ _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14708__I _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11867_ _06774_ register_file\[6\]\[3\] _06775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13612__I _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15770__CLK clknet_leaf_255_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08068__A1 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13606_ _01121_ _01124_ _01126_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_158_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10818_ _06095_ _06096_ _06097_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08706__I _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14586_ _01110_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09804__A2 register_file\[21\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11798_ _06660_ _06730_ _06733_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16325_ _00713_ clknet_leaf_77_clk register_file\[20\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12228__I _06090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13537_ _00998_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11611__A2 _06602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10749_ _06040_ _06041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_158_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16126__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16256_ _00644_ clknet_5_3__leaf_clk register_file\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13468_ _07578_ _07730_ _07772_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13768__B _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09568__A1 _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15207_ _02707_ _02709_ _02544_ _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12419_ _07009_ _07112_ _07118_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16187_ _00575_ clknet_leaf_40_clk register_file\[25\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11375__A1 _06462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13399_ _07509_ _07728_ _07732_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15138_ _02474_ register_file\[16\]\[18\] _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10192__B _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15069_ _02569_ _02572_ _02242_ _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07960_ _01175_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11127__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_4_clk clknet_5_0__leaf_clk clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12875__A1 _07359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07891_ _01062_ _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09630_ _04936_ _04941_ _04002_ _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09740__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10350__A2 register_file\[18\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14616__A2 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09561_ _04869_ _04872_ _04873_ _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12627__A1 _07244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08512_ _03826_ _03834_ _03838_ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09492_ _04804_ _04805_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10102__A2 register_file\[22\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08443_ _03769_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11850__A2 _06758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13522__I _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08374_ _03701_ register_file\[8\]\[31\] _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08059__A1 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13052__A1 _07511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07806__A1 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11602__A2 _06602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_18__f_clk clknet_3_4_0_clk clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10169__A2 register_file\[24\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11366__A1 _06388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08782__A2 register_file\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11118__A1 _06108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15643__CLK clknet_leaf_271_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11669__A2 register_file\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12866__A1 _07295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15184__I _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09828_ _05002_ register_file\[9\]\[18\] _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14607__A2 register_file\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09759_ _05065_ _05068_ _04102_ _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08298__A1 _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12770_ _07340_ register_file\[20\]\[19\] _07342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12094__A2 _06866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11721_ _06675_ register_file\[8\]\[15\] _06681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13432__I _07737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16149__CLK clknet_leaf_181_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14440_ _01951_ _01786_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11652_ _06434_ _06630_ _06632_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10603_ _03821_ register_file\[9\]\[30\] _05900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14371_ _01882_ _01883_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11583_ _06024_ _04001_ _06590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16110_ _00498_ clknet_leaf_192_clk register_file\[3\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13322_ _07681_ _07686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10534_ _05637_ register_file\[2\]\[28\] _05833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16299__CLK clknet_leaf_138_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13346__A2 _07697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16041_ _00429_ clknet_leaf_291_clk register_file\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13253_ _07638_ register_file\[14\]\[7\] _07645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10465_ _05755_ _05764_ _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11357__A1 _06454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12204_ _06059_ _06980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13184_ _07534_ _07601_ _07603_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10396_ _05694_ _05696_ _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15099__A2 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12135_ _06677_ _06929_ _06935_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08773__A2 register_file\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14846__A2 _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12857__A1 _07388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12066_ _06892_ net21 _06894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11017_ _06073_ _06236_ _06237_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10332__A2 register_file\[31\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15825_ _00213_ clknet_leaf_170_clk register_file\[26\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14074__A3 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15756_ _00144_ clknet_leaf_136_clk register_file\[13\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08289__A1 _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13282__A1 _07660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12968_ _07458_ register_file\[17\]\[2\] _07461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10096__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14707_ _02045_ _02213_ _02215_ _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11919_ _06701_ _06799_ _06805_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15687_ _00075_ clknet_leaf_85_clk register_file\[28\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11832__A2 _06751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12899_ _07414_ register_file\[18\]\[6\] _07420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14638_ _01980_ register_file\[26\]\[12\] _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13034__A1 _07304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14882__B _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09789__A1 _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13585__A2 _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14569_ _02078_ _01914_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11596__A1 _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10399__A2 register_file\[9\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16308_ _00696_ clknet_leaf_180_clk register_file\[21\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08090_ _03419_ _01141_ _03421_ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16239_ _00627_ clknet_leaf_153_clk register_file\[23\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13337__A2 _07690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14173__I _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11348__A1 _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15666__CLK clknet_leaf_178_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08213__A1 _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08992_ _04029_ register_file\[17\]\[6\] _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14837__A2 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07943_ _03276_ register_file\[15\]\[25\] _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12848__A1 _07388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09713__A1 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07874_ _03202_ _03208_ _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10323__A2 register_file\[26\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09613_ _04921_ _04924_ _04452_ _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09544_ _04854_ _04856_ _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13273__A1 _07653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12076__A2 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09475_ _04516_ register_file\[26\]\[13\] _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08426_ _03706_ register_file\[20\]\[31\] _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13025__A1 _07491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08357_ _03682_ _03684_ _01045_ _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ _03613_ _03616_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11339__A1 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10250_ _05551_ _05552_ _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16591__CLK clknet_leaf_189_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10011__A1 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14811__I _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10181_ _05482_ _05484_ _05485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10116__I _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14828__A2 register_file\[18\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12839__A1 _07269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13427__I _07729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14032__B _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13940_ _01177_ _01453_ _01457_ _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_59_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09126__B _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11511__A1 _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13871_ _01039_ register_file\[21\]\[3\] _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08965__B _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15610_ _01074_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12822_ _07252_ _07370_ _07373_ _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13264__A1 _07534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16590_ _00978_ clknet_leaf_188_clk register_file\[9\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12067__A2 _06888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10078__A1 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15541_ register_file\[4\]\[22\] _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12753_ _07326_ register_file\[20\]\[12\] _07332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10786__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11814__A2 register_file\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13162__I _07585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11704_ _06663_ register_file\[8\]\[10\] _06669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13016__A1 _07286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15472_ _02963_ _02971_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12684_ _06121_ _07286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14423_ _01933_ _01934_ _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11635_ _06417_ _06616_ _06622_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13567__A2 _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11578__A1 _06440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14354_ _01865_ _01694_ _01866_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11566_ _06579_ register_file\[11\]\[24\] _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15089__I _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13305_ _07631_ register_file\[14\]\[29\] _07675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13319__A2 _07680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10517_ _05814_ _05815_ _05816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14285_ _01623_ _01796_ _01798_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_155_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11497_ _06495_ register_file\[12\]\[29\] _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09087__I _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16024_ _00412_ clknet_leaf_243_clk register_file\[6\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13236_ _07634_ register_file\[14\]\[0\] _07635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10448_ _05483_ register_file\[4\]\[27\] _05748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08746__A2 register_file\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10026__I _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13167_ _07585_ _07593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10379_ _05676_ _05679_ _04078_ _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10553__A2 register_file\[19\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12118_ _06660_ _06922_ _06925_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13098_ _07543_ _07544_ _07545_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12241__I _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12049_ _06878_ net14 _06884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11502__A1 _06444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14877__B _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09171__A2 register_file\[12\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15552__I _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15808_ _00196_ clknet_leaf_10_clk register_file\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12058__A2 _06888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10069__A1 _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15739_ _00127_ clknet_5_7__leaf_clk register_file\[27\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16464__CLK clknet_leaf_166_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13072__I _07506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09260_ _04576_ register_file\[31\]\[10\] _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08211_ _03540_ _02978_ _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09191_ _04441_ register_file\[14\]\[9\] _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13800__I _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11569__A1 _06579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08142_ _03469_ _03472_ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12230__A2 _06988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14507__A1 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08073_ _03401_ _03404_ _03075_ _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08985__A2 register_file\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_295_clk clknet_5_4__leaf_clk clknet_leaf_295_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15180__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11741__A1 _06687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08975_ _04280_ _04296_ _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13247__I _07633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07926_ _03252_ _03259_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12297__A2 _07040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input25_I new_value[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09162__A2 register_file\[24\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07857_ _03027_ register_file\[13\]\[24\] _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15235__A2 register_file\[22\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12049__A2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13246__A1 _07516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07788_ _02786_ _03123_ _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09527_ _04840_ _04637_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14994__A1 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09458_ _04633_ register_file\[1\]\[12\] _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08673__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08409_ _03736_ _03657_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09389_ _04633_ register_file\[1\]\[11\] _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11420_ _06442_ _06450_ _06492_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10555__B _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14027__B _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_286_clk clknet_5_5__leaf_clk clknet_leaf_286_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10232__A1 _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11351_ _06373_ _06448_ _06452_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output93_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11980__A1 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10302_ _05338_ register_file\[13\]\[25\] _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15171__A1 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14070_ _01327_ register_file\[23\]\[5\] _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11282_ _06403_ register_file\[19\]\[13\] _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13021_ _07290_ _07487_ _07492_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09925__A1 _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13721__A2 register_file\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10233_ _05334_ register_file\[11\]\[24\] _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11732__A1 _06686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10535__A2 register_file\[3\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16337__CLK clknet_leaf_157_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10164_ _05332_ register_file\[10\]\[23\] _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14972_ _02475_ _02476_ _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10095_ _05332_ register_file\[30\]\[22\] _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_clk_I clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10299__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09153__A2 register_file\[9\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13923_ _01433_ _01440_ _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16487__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15226__A2 register_file\[19\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_210_clk clknet_5_23__leaf_clk clknet_leaf_210_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08900__A2 register_file\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13237__A1 _07502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13854_ _01368_ _01372_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12805_ _07230_ _07360_ _07363_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16573_ _00961_ clknet_leaf_304_clk register_file\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13785_ _01300_ _01303_ _01052_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10997_ _06220_ _06225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15524_ _03021_ _03022_ _02691_ _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12736_ _07321_ _07322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12460__A2 _07136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14737__A1 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15455_ register_file\[4\]\[21\] _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12667_ _06099_ _07274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13620__I _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14406_ _01835_ register_file\[18\]\[9\] _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11618_ _06400_ _06609_ _06612_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12212__A2 register_file\[31\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15386_ _02864_ _02885_ _02886_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12598_ _07028_ _07222_ _07225_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10223__A1 _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_277_clk clknet_5_7__leaf_clk clknet_leaf_277_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14337_ _01508_ register_file\[8\]\[8\] _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08967__A2 register_file\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11549_ _06565_ register_file\[11\]\[17\] _06571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13960__A2 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10774__A2 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14268_ _01778_ _01781_ _01608_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_171_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09916__A1 _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16007_ _00395_ clknet_leaf_297_clk register_file\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13219_ _07619_ register_file\[15\]\[26\] _07624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13712__A2 register_file\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14199_ _01713_ register_file\[2\]\[6\] _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10526__A2 _05824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15465__A2 register_file\[2\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14268__A3 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15704__CLK clknet_leaf_196_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08760_ _04079_ _04084_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12279__A2 register_file\[31\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09144__A2 register_file\[20\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08691_ _04014_ _04015_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_201_clk clknet_5_19__leaf_clk clknet_leaf_201_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13228__A1 _07578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15854__CLK clknet_leaf_126_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14976__A1 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11315__I _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09312_ _04625_ _04628_ _04002_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14728__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09243_ _04492_ register_file\[30\]\[9\] _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10462__A1 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13530__I _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08407__A1 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09174_ _04492_ register_file\[14\]\[8\] _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12203__A2 _06976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13400__A1 _07730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08958__A2 _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08125_ _03456_ _03132_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11962__A1 _06830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15153__A1 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08056_ _03365_ _03388_ _03303_ _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_150_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15457__I register_file\[5\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14900__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput49 net49 rD[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11714__A1 _06675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09383__A2 register_file\[18\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11190__A2 register_file\[13\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08958_ _04272_ _04279_ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13467__A1 _07727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07909_ _01107_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08889_ _04211_ register_file\[13\]\[4\] _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13705__I _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10920_ _06177_ _06178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13219__A1 _07619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08894__A1 _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10851_ net25 _06124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13570_ _01090_ register_file\[30\]\[0\] _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10782_ _06067_ _06068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12442__A2 _07126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12521_ _07135_ register_file\[23\]\[29\] _07179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10453__A1 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08110__A3 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15240_ _02731_ _02741_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12452_ _07138_ register_file\[23\]\[0\] _07139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08534__I _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10205__A1 _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11403_ _06446_ _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_259_clk clknet_5_19__leaf_clk clknet_leaf_259_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_184_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15171_ _02673_ register_file\[29\]\[18\] _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12056__I _06873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12383_ _07089_ _07097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09071__A1 _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11953__A1 _06822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10756__A2 register_file\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14122_ _01550_ register_file\[25\]\[6\] _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15144__A1 _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11334_ _06155_ _06440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15727__CLK clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14053_ _01567_ _01480_ _01568_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14271__I register_file\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11265_ _06391_ register_file\[19\]\[8\] _06392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11705__A1 _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13004_ _07274_ _07480_ _07482_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10216_ _05248_ register_file\[19\]\[24\] _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09374__A2 register_file\[10\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11196_ _06100_ _06344_ _06346_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11181__A2 register_file\[13\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15447__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10147_ _05448_ _05450_ _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13458__A1 _07567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14955_ _02460_ _02378_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10078_ _05117_ register_file\[18\]\[22\] _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12130__A1 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14670__A3 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13906_ _01423_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14886_ _02389_ _02391_ _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13837_ _01353_ _01355_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10692__A1 _05980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16556_ _00944_ clknet_leaf_130_clk register_file\[29\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13768_ _01240_ _01287_ _01201_ net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15507_ _03004_ _02672_ _03005_ _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12719_ _06216_ _03836_ _07310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16487_ _00875_ clknet_leaf_48_clk register_file\[15\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_0_clk clk clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13699_ _01214_ _01218_ _01052_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15438_ _02935_ _02937_ _02691_ _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14186__A2 _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_274_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07860__A2 register_file\[15\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15369_ register_file\[4\]\[20\] _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11944__A1 _06818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15135__A1 _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_289_clk_I clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09930_ _05173_ register_file\[3\]\[19\] _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13697__A1 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08168__A3 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09861_ _05167_ _05169_ _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11172__A2 _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ _03986_ register_file\[30\]\[3\] _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_212_clk_I clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09792_ _04832_ register_file\[15\]\[17\] _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13449__A1 _07756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09117__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08743_ _04067_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14110__A2 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12121__A1 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13525__I _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08876__A1 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ _03998_ _03999_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12672__A2 _07272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16032__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_4__f_clk_I clknet_3_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08628__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12424__A2 _07119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10435__A1 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13260__I _07641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10986__A2 _06216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09226_ _04409_ register_file\[11\]\[9\] _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14177__A2 register_file\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07851__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12188__A1 _06967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09157_ _04407_ register_file\[10\]\[8\] _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09053__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13924__A2 register_file\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11935__A1 _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15126__A1 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08108_ _03276_ register_file\[15\]\[27\] _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09088_ _04407_ register_file\[10\]\[7\] _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ _03203_ _03371_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13688__A1 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09356__A2 register_file\[30\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11050_ _06135_ _06250_ _06256_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12360__A1 _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11163__A2 register_file\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10001_ _05304_ _05305_ _05307_ _05308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09108__A2 register_file\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output56_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14740_ _02247_ _01914_ _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09134__B _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11952_ _06825_ _06826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_40_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13860__A1 _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10903_ _06024_ _04636_ _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10674__A1 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14671_ _02168_ _02179_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08331__A3 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11883_ _06665_ _06778_ _06784_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16410_ _00798_ clknet_leaf_272_clk register_file\[18\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13622_ _01142_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15601__A2 register_file\[8\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10834_ _06108_ _06096_ _06110_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08619__A1 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16525__CLK clknet_leaf_125_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16341_ _00729_ clknet_leaf_206_clk register_file\[20\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10794__I _06077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13553_ _01024_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_41_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09292__A1 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10765_ net39 _06054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08095__A2 register_file\[9\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12504_ _07014_ _07167_ _07169_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16272_ _00660_ clknet_leaf_155_clk register_file\[22\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14168__A2 register_file\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15365__A1 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13484_ _01004_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10696_ _05990_ _05991_ _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15223_ _02723_ _02724_ _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12435_ _07123_ register_file\[24\]\[26\] _07128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13915__A2 _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11926__A1 _06708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15154_ _02655_ _02323_ _02656_ _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_148_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12366_ _07036_ _07042_ _07085_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14105_ _01615_ _01620_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11317_ _06426_ _06420_ _06428_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15085_ _02587_ _02257_ _02588_ _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12297_ _06967_ _07040_ _07045_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14036_ _01549_ _01551_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11248_ _06377_ _06369_ _06379_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12351__A1 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10034__I _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11179_ _06069_ _06330_ _06336_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15987_ _00375_ clknet_leaf_228_clk register_file\[7\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12103__A1 _06645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08439__I _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14938_ _01455_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08858__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12654__A2 register_file\[21\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10665__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14869_ _02373_ _02375_ _02127_ _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12406__A2 register_file\[24\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08390_ _03716_ _01046_ _03717_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13603__A1 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10417__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08086__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16539_ _00927_ clknet_leaf_287_clk register_file\[14\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11090__A1 _06275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_93_clk_I clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09011_ _04330_ _04331_ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09035__A1 _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11917__A1 _06698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11393__A2 _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12590__A1 _07219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09219__B _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ _05090_ register_file\[20\]\[19\] _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14331__A2 register_file\[22\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_151_clk_I clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12342__A1 _07011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11145__A2 _06271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09844_ _05151_ _05152_ _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12893__A2 register_file\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09775_ _05084_ register_file\[7\]\[17\] _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10879__I _06146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13255__I _07633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_166_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08726_ _04049_ _04050_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12645__A2 _07248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16548__CLK clknet_leaf_69_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14795__B _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10656__A1 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08657_ _03880_ register_file\[21\]\[1\] _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_46_clk_I clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15595__A1 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08588_ _03903_ _03910_ _03914_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_168_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10408__A1 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09274__A1 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13070__A2 _07520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10959__A2 register_file\[2\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11081__A1 _06041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10550_ _05589_ register_file\[16\]\[29\] _05848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09209_ _04320_ register_file\[7\]\[9\] _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_104_clk_I clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09026__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14814__I _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10481_ _03821_ register_file\[17\]\[28\] _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12220_ _06990_ _06988_ _06991_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14570__A2 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10563__B _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12581__A1 _07212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12151_ _06940_ register_file\[3\]\[21\] _06945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11102_ _06283_ register_file\[27\]\[12\] _06289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12082_ _03287_ _06902_ _06903_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12333__A1 _07061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11136__A2 register_file\[27\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11033_ _06104_ _06243_ _06246_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15910_ _00298_ clknet_leaf_109_clk register_file\[10\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08001__A2 register_file\[28\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10789__I _06051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15841_ _00229_ clknet_leaf_22_clk register_file\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12984_ _07470_ register_file\[17\]\[8\] _07471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15772_ _00160_ clknet_leaf_279_clk register_file\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13833__A1 _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10647__A1 _05940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14723_ _02230_ register_file\[27\]\[13\] _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11935_ _06317_ _03912_ _06814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15915__CLK clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14654_ _02162_ _01832_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11866_ _06769_ _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13605_ _01125_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10817_ _06087_ register_file\[30\]\[15\] _06097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14585_ _01932_ register_file\[8\]\[11\] _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11797_ _06726_ register_file\[7\]\[7\] _06733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16324_ _00712_ clknet_leaf_73_clk register_file\[20\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15338__A1 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13536_ _01056_ register_file\[24\]\[0\] _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10748_ _06039_ _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16255_ _00643_ clknet_leaf_24_clk register_file\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13467_ _07727_ register_file\[9\]\[30\] _07772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10679_ _05731_ register_file\[28\]\[31\] _05975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15206_ _02708_ _02542_ _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12418_ _07116_ register_file\[24\]\[19\] _07118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16186_ _00574_ clknet_leaf_40_clk register_file\[25\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13398_ _07730_ register_file\[9\]\[1\] _07732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12572__A1 _07002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15137_ _02598_ _02640_ _02473_ net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12349_ _07018_ _07071_ _07076_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15068_ _02570_ _02323_ _02571_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12324__A1 _07061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11127__A2 _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14019_ _01533_ _01535_ _01273_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07890_ _03221_ _03223_ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12875__A2 register_file\[1\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10886__A1 _06026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13075__I _06067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09560_ _04219_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_110_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12627__A2 _07233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08511_ _03837_ _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10638__A1 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09491_ _04602_ register_file\[23\]\[13\] _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08442_ net1 net2 _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09256__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08373_ _01179_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_17_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13052__A2 _07505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11063__A1 _06160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07806__A2 register_file\[17\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14001__A1 _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08632__I _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14552__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11366__A2 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15501__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12315__A1 _06985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11118__A2 _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12866__A2 _07398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16370__CLK clknet_leaf_159_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09827_ _05132_ _05135_ _03877_ _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10877__A1 _06144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15938__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _05066_ _05067_ _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13815__A1 _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08709_ _03956_ register_file\[10\]\[2\] _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10629__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09689_ _04997_ _04999_ _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08298__A2 register_file\[25\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11720_ _06655_ _06680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08807__I _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11651_ _06627_ register_file\[10\]\[26\] _06632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09247__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11233__I _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11054__A1 _06254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10602_ _05870_ _05899_ _05647_ net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14370_ _01155_ _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11582_ _06444_ _06546_ _06589_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13321_ _07511_ _07680_ _07685_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10801__A1 _06082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10533_ _05828_ _05831_ _05028_ _05832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_195_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16040_ _00428_ clknet_leaf_296_clk register_file\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13252_ _07522_ _07642_ _07644_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10464_ _05760_ _05763_ _03816_ _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10293__B _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12554__A1 _07198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12203_ _06978_ _06976_ _06979_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13183_ _07598_ register_file\[15\]\[11\] _07603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10395_ _05695_ register_file\[23\]\[26\] _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12134_ _06933_ register_file\[3\]\[14\] _06935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12306__A1 _06974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12065_ _02706_ _06888_ _06893_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12857__A2 register_file\[1\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09373__I _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11016_ _06233_ register_file\[28\]\[10\] _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11408__I _06457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15824_ _00212_ clknet_leaf_169_clk register_file\[26\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_24__f_clk clknet_3_6_0_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15755_ _00143_ clknet_leaf_136_clk register_file\[13\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12967_ _07237_ _07456_ _07460_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11293__A1 _06410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14706_ _02214_ _01883_ _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10096__A2 register_file\[31\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11918_ _06803_ register_file\[6\]\[24\] _06805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15559__A1 _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15686_ _00074_ clknet_leaf_83_clk register_file\[28\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12898_ _07246_ _07418_ _07419_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14637_ _01813_ register_file\[27\]\[12\] _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11849_ _06719_ register_file\[7\]\[29\] _06763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13034__A2 _07494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11045__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14568_ _02076_ _02077_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13585__A3 _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12793__A1 _07311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11596__A2 _06592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16307_ _00695_ clknet_leaf_209_clk register_file\[21\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16243__CLK clknet_leaf_181_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13519_ _01039_ register_file\[21\]\[0\] _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14499_ _02006_ _02009_ _01671_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_146_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16238_ _00626_ clknet_leaf_145_clk register_file\[23\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12545__A1 _07190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11348__A2 register_file\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16169_ _00557_ clknet_leaf_93_clk register_file\[25\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09410__A1 _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08213__A2 register_file\[18\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16393__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08991_ _04304_ _04311_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15285__I register_file\[4\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07972__A1 _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07942_ _01455_ _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12848__A2 register_file\[1\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09283__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07873_ _03205_ _03207_ _02960_ _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11318__I _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ _04922_ _04923_ _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10222__I _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09543_ _04855_ register_file\[27\]\[14\] _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14470__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13273__A2 register_file\[14\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09474_ _04786_ _04787_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08425_ _03750_ _03752_ _01159_ _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09229__A1 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14222__A1 _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11036__A1 _06108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08356_ _03683_ _01059_ _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14773__A2 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11988__I _06825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08287_ _03614_ _03615_ _01076_ _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_192_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14525__A2 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12536__A1 _07186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11339__A2 _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09401__A1 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10011__A2 register_file\[22\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10180_ _05483_ register_file\[4\]\[23\] _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15760__CLK clknet_leaf_173_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12612__I _07234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12839__A2 _07377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11511__A2 _06544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13870_ _01387_ register_file\[20\]\[3\] _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16116__CLK clknet_leaf_221_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12821_ _07366_ register_file\[1\]\[7\] _07373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__A1 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14461__A1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13264__A2 _07649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12752_ _07262_ _07329_ _07331_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10078__A2 register_file\[18\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11275__A1 _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15540_ _03035_ _03038_ _02953_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09142__B _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08537__I _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08140__A1 _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11703_ _06655_ _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_37_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15471_ _02970_ _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16266__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12683_ _07283_ _07284_ _07285_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13016__A2 _07487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14213__A1 _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14422_ _01676_ register_file\[9\]\[9\] _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11634_ _06620_ register_file\[10\]\[19\] _06622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12775__A1 _07340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11578__A2 _06582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14353_ _01605_ register_file\[15\]\[8\] _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11565_ _06426_ _06575_ _06580_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09640__A1 _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13304_ _07574_ _07670_ _07674_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10516_ _05752_ register_file\[11\]\[28\] _05815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14284_ _01797_ _01456_ _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11496_ _06438_ _06534_ _06538_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16023_ _00411_ clknet_5_20__leaf_clk register_file\[6\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13235_ _07633_ _07634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_155_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10447_ _05481_ register_file\[5\]\[27\] _05747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10307__I _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13166_ _07516_ _07584_ _07592_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ _05677_ _05678_ _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07954__A1 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13618__I _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14819__A3 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12117_ _06918_ register_file\[3\]\[7\] _06925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13097_ _07539_ register_file\[16\]\[15\] _07545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12048_ _02122_ _06881_ _06883_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11502__A2 _06498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15807_ _00195_ clknet_leaf_11_clk register_file\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14449__I _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13999_ _01514_ _01515_ _01431_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11266__A1 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10069__A2 register_file\[1\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15738_ _00126_ clknet_leaf_267_clk register_file\[27\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09987__B _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15669_ _00057_ clknet_leaf_224_clk register_file\[2\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08682__A2 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08210_ _03539_ _03225_ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11018__A1 _06233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09190_ _04506_ _04507_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14755__A2 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15633__CLK clknet_leaf_165_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12766__A1 _07276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11569__A2 register_file\[11\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08141_ _03470_ _03471_ _03231_ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08434__A2 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08072_ _03402_ _03155_ _03403_ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12518__A1 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13191__A1 _07541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11741__A2 register_file\[8\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12432__I _07097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08974_ _04287_ _04295_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16139__CLK clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07925_ _03255_ _03258_ _02924_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07856_ _02940_ register_file\[12\]\[24\] _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input18_I new_value[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07787_ register_file\[4\]\[23\] _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13246__A2 _07632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09526_ _04836_ _04838_ _04839_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14994__A2 register_file\[18\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09457_ _04499_ register_file\[3\]\[12\] _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11009__A1 _06060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08408_ register_file\[27\]\[31\] _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09388_ _04499_ register_file\[3\]\[11\] _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12757__A1 _07266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08339_ register_file\[5\]\[30\] _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12607__I _06020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09622__A1 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11350_ _06450_ register_file\[26\]\[1\] _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12509__A1 _07018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10301_ _05599_ _05602_ _05268_ _05603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11980__A2 _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11281_ _06370_ _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13020_ _07491_ register_file\[17\]\[23\] _07492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13182__A1 _07531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output86_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10232_ _05332_ register_file\[10\]\[24\] _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09925__A2 register_file\[10\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11732__A2 _06680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10163_ _05465_ _05466_ _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14971_ _02390_ register_file\[25\]\[16\] _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10094_ _05396_ _05398_ _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14682__A1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13922_ _01436_ _01439_ _01148_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11496__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10299__A2 register_file\[11\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10797__I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13853_ _01369_ register_file\[1\]\[2\] _01371_ _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14434__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13237__A2 _07632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12804_ _07362_ register_file\[1\]\[0\] _07363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11248__A1 _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16572_ _00960_ clknet_leaf_286_clk register_file\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15656__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14985__A2 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13784_ _01301_ _01046_ _01302_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10996_ _06037_ _06219_ _06224_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12996__A1 _07477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15523_ _02936_ register_file\[10\]\[22\] _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12735_ _07313_ _07321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12666_ _07271_ _07272_ _07273_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15454_ _02950_ _02952_ _02953_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14405_ _01746_ register_file\[19\]\[9\] _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11617_ _06606_ register_file\[10\]\[12\] _06612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12597_ _07219_ register_file\[22\]\[27\] _07225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15385_ _01193_ _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11420__A1 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14336_ _01827_ _01848_ _01506_ _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11548_ _06410_ _06568_ _06570_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14267_ _01779_ _01694_ _01780_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15162__A2 _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11479_ _06524_ register_file\[12\]\[21\] _06529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13173__A1 _07590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16006_ _00394_ clknet_leaf_309_clk register_file\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13218_ _07567_ _07622_ _07623_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09916__A2 register_file\[23\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14198_ _01277_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_140_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12252__I _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13149_ _07504_ register_file\[16\]\[31\] _07581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14673__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08886__B _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16431__CLK clknet_leaf_144_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11487__A1 _06429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08690_ _03786_ register_file\[19\]\[2\] _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14179__I _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13228__A2 _07586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09311_ _04626_ _04627_ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12987__A1 _07257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09242_ _04557_ _04559_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10462__A2 register_file\[31\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12739__A1 _07318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14128__B _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12427__I _07086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09173_ _04145_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13400__A2 register_file\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11331__I _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08124_ register_file\[3\]\[27\] _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11411__A1 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11962__A2 register_file\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08055_ _03379_ _03387_ _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15153__A2 register_file\[23\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07965__B _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13164__A1 _07513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12911__A1 _07422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11714__A2 register_file\[8\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08591__A1 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08957_ _04275_ _04278_ _04068_ _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13467__A2 register_file\[9\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11478__A1 _06419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07908_ _03233_ _03241_ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08888_ _03897_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15679__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08343__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14089__I _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07839_ _03007_ register_file\[30\]\[24\] _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10150__A1 _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13219__A2 register_file\[15\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11506__I _06542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10850_ _06122_ _06118_ _06123_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12978__A1 _07246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ _04691_ register_file\[31\]\[13\] _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10781_ net42 _06067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09843__A1 _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12520_ _07030_ _07174_ _07178_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09420__B _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11650__A1 _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14719__A2 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08815__I _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12451_ _07137_ _07138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_166_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14195__A3 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11402_ _06424_ _06479_ _06482_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11402__A1 _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15170_ _01134_ _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10205__A2 register_file\[3\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16304__CLK clknet_leaf_158_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12382_ _06972_ _07088_ _07096_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09071__A2 register_file\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14121_ _01635_ register_file\[24\]\[6\] _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11953__A2 register_file\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11333_ _06438_ _06432_ _06439_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_21__f_clk_I clknet_3_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14052_ _01216_ register_file\[31\]\[5\] _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11264_ _06370_ _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08550__I _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13003_ _07477_ register_file\[17\]\[16\] _07482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12902__A1 _07252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13168__I _07593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11705__A2 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10215_ _05452_ register_file\[18\]\[24\] _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11195_ _06341_ register_file\[13\]\[16\] _06346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08582__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10146_ _05449_ register_file\[28\]\[23\] _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13458__A2 _07766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11469__A1 _06517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12800__I _07358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ _05380_ _05381_ _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14954_ _02454_ _02459_ _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12130__A2 _06929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13905_ _01004_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14885_ _02390_ register_file\[25\]\[15\] _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_195_clk clknet_5_18__leaf_clk clknet_leaf_195_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13836_ _01354_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12969__A1 _07239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14727__I _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16555_ _00943_ clknet_leaf_134_clk register_file\[29\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08637__A2 _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13767_ _01262_ _01286_ _01195_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10979_ _06167_ register_file\[2\]\[30\] _06212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13631__I _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15506_ _02673_ register_file\[29\]\[22\] _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11641__A1 _06620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12718_ _07308_ _07235_ _07309_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16486_ _00874_ clknet_leaf_48_clk register_file\[15\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13698_ _01215_ _01046_ _01217_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15437_ _02936_ register_file\[10\]\[21\] _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12649_ _07259_ _07260_ _07261_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15368_ _02866_ _02868_ _02537_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14462__I _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14319_ _01009_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10990__I _06220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15299_ _02800_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13146__A1 _07504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13697__A2 register_file\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09860_ _05168_ register_file\[27\]\[18\] _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08811_ _04133_ _04134_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09791_ _04830_ register_file\[14\]\[17\] _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13449__A2 register_file\[9\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13806__I _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08742_ _03794_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12710__I _06155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08325__A1 _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12121__A2 _06922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08673_ _03908_ register_file\[11\]\[1\] _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_186_clk clknet_5_28__leaf_clk clknet_leaf_186_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10132__A1 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15971__CLK clknet_leaf_314_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11880__A1 _06782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15071__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09825__A1 _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08628__A2 register_file\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13541__I _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11632__A1 _06620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10435__A2 register_file\[11\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16327__CLK clknet_leaf_80_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09225_ _04407_ register_file\[10\]\[9\] _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12188__A2 _06961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13385__A1 _07679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09156_ _04472_ _04474_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_5_clk_I clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08107_ _03274_ register_file\[14\]\[27\] _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16477__CLK clknet_leaf_301_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15126__A2 register_file\[2\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09087_ _03867_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_clk clknet_5_13__leaf_clk clknet_leaf_110_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_107_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13137__A1 _07563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08038_ register_file\[4\]\[26\] _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_190_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14885__A1 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10000_ _05306_ register_file\[1\]\[20\] _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08564__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12360__A2 _07078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09989_ _05228_ register_file\[21\]\[20\] _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14637__A1 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_5__f_clk clknet_3_1_0_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08316__A1 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output49_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10123__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_177_clk clknet_5_29__leaf_clk clknet_leaf_177_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11951_ _06817_ _06825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_177_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11236__I _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13860__A2 register_file\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10902_ _06164_ _06029_ _06165_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14670_ _02172_ _02178_ _02091_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11882_ _06782_ register_file\[6\]\[9\] _06784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10674__A2 register_file\[23\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10833_ _06109_ register_file\[30\]\[18\] _06110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13621_ _01095_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14547__I _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09816__A1 _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13451__I _07726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11623__A1 _06405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16340_ _00728_ clknet_leaf_180_clk register_file\[20\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10764_ _06050_ _06052_ _06053_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13552_ _01072_ register_file\[26\]\[0\] _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09292__A2 register_file\[12\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12503_ _07164_ register_file\[23\]\[21\] _07169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16271_ _00659_ clknet_leaf_154_clk register_file\[22\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13483_ _01003_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15365__A2 register_file\[6\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10695_ _03844_ register_file\[4\]\[31\] _05991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07842__A3 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15222_ _02390_ register_file\[17\]\[19\] _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12434_ _07023_ _07126_ _07127_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15378__I register_file\[3\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11926__A2 _06806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15153_ _02488_ register_file\[23\]\[18\] _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12365_ _07039_ register_file\[25\]\[31\] _07085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15117__A2 _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_101_clk clknet_5_15__leaf_clk clknet_leaf_101_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_165_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13128__A1 _07565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11316_ _06427_ register_file\[19\]\[23\] _06428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14104_ _01617_ _01619_ _01273_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_153_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15084_ _02258_ register_file\[21\]\[17\] _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15844__CLK clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12296_ _07042_ register_file\[25\]\[2\] _07045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14876__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14035_ _01550_ register_file\[25\]\[5\] _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11247_ _06378_ register_file\[19\]\[3\] _06379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12351__A2 _07071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11178_ _06334_ register_file\[13\]\[9\] _06336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10362__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13626__I _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15994__CLK clknet_leaf_252_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10129_ _05230_ register_file\[8\]\[22\] _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12530__I _07182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09325__B _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15986_ _00374_ clknet_leaf_229_clk register_file\[7\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08307__A1 _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12103__A2 _06912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13300__A1 _07570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14937_ _02442_ register_file\[14\]\[15\] _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10114__A1 _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_168_clk clknet_5_31__leaf_clk clknet_leaf_168_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11862__A1 _06770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10665__A2 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14868_ _02374_ _02125_ _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15053__A1 _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13819_ _01247_ register_file\[11\]\[2\] _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14799_ _02286_ _02306_ _02054_ _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14800__A1 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11614__A1 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16538_ _00926_ clknet_leaf_254_clk register_file\[14\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09995__B _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11090__A2 register_file\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14159__A3 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16469_ _00857_ clknet_leaf_215_clk register_file\[16\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09010_ _04259_ register_file\[23\]\[6\] _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13367__A1 _07708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09035__A2 register_file\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11917__A2 _06799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14192__I _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15108__A2 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08190__I register_file\[4\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09912_ _05088_ register_file\[21\]\[19\] _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12342__A2 _07071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09843_ _05084_ register_file\[31\]\[18\] _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08010__A3 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09774_ _03850_ _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08725_ _03864_ register_file\[4\]\[2\] _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_159_clk clknet_5_31__leaf_clk clknet_leaf_159_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13842__A2 _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11853__A1 _06719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10656__A2 register_file\[2\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08656_ _03978_ _03981_ _03877_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15044__A1 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10895__I _06159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08587_ _03913_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15717__CLK clknet_leaf_69_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11605__A1 _06598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10408__A2 register_file\[1\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15347__A2 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11081__A2 _06269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13358__A1 _07548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09208_ _04317_ register_file\[6\]\[9\] _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10480_ _05746_ _05779_ _05647_ net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09139_ _04317_ register_file\[6\]\[8\] _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12615__I _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08785__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12581__A2 register_file\[22\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12150_ _06691_ _06943_ _06944_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10592__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11101_ _06078_ _06286_ _06288_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12081_ _06899_ net28 _06903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12333__A2 register_file\[25\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11032_ _06240_ register_file\[28\]\[17\] _06246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15840_ _00228_ clknet_leaf_5_clk register_file\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14086__A2 _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15771_ _00159_ clknet_leaf_283_clk register_file\[13\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12983_ _07457_ _07470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14722_ _01014_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11844__A1 _06706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11934_ _06716_ _06770_ _06813_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15035__A1 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14653_ _02161_ _01914_ _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14277__I register_file\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_288_clk_I clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11865_ _06647_ _06768_ _06773_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13604_ _01074_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10816_ _06051_ _06096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14584_ _02075_ _02093_ _01930_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11796_ _06658_ _06730_ _06732_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16323_ _00711_ clknet_leaf_68_clk register_file\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13535_ _01055_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15338__A2 register_file\[22\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10747_ net36 _06039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_211_clk_I clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13349__A1 _07538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16254_ _00642_ clknet_leaf_43_clk register_file\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13466_ _07576_ _07766_ _07771_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10678_ _05729_ register_file\[29\]\[31\] _05974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15205_ register_file\[5\]\[18\] _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12417_ _07006_ _07112_ _07117_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16185_ _00573_ clknet_leaf_196_clk register_file\[25\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13397_ _07502_ _07728_ _07731_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08776__A1 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12572__A2 _07208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15136_ _02617_ _02639_ _02471_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12348_ _07075_ register_file\[25\]\[23\] _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10583__A1 _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_226_clk_I clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14849__A1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15067_ _02488_ register_file\[31\]\[17\] _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12279_ _06960_ register_file\[31\]\[29\] _07033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14313__A3 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12324__A2 register_file\[25\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14018_ _01534_ _01271_ _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09055__B _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16172__CLK clknet_leaf_138_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15969_ _00357_ clknet_leaf_314_clk register_file\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08510_ _03836_ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09490_ _04600_ register_file\[22\]\[13\] _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08441_ _03767_ register_file\[25\]\[0\] _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14187__I _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13588__A1 _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08372_ _03699_ _01011_ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09256__A2 register_file\[28\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12260__A1 _07019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15329__A2 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11063__A2 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_313_clk clknet_5_0__leaf_clk clknet_leaf_313_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_176_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12012__A1 _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08767__A1 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10574__A1 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14650__I _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12315__A2 _07050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16515__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10326__A1 _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09192__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09826_ _05133_ _05134_ _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10877__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14068__A2 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12079__A1 _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09757_ _04998_ register_file\[19\]\[17\] _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13815__A2 register_file\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11826__A1 _06748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08708_ _04030_ _04032_ _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10629__A2 register_file\[19\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09688_ _04998_ register_file\[7\]\[16\] _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ _03964_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14097__I register_file\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11514__I _06545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11650_ _06431_ _06630_ _06631_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09247__A2 register_file\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14240__A2 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10601_ _05885_ _05898_ _05899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12251__A1 _07011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11054__A2 register_file\[28\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11581_ _06543_ register_file\[11\]\[31\] _06589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_304_clk clknet_5_1__leaf_clk clknet_leaf_304_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_22_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13320_ _07682_ register_file\[29\]\[2\] _07685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10532_ _05829_ _05830_ _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10801__A2 _06074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12003__A1 _06851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10463_ _05761_ _05762_ _05763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13251_ _07638_ register_file\[14\]\[6\] _07644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12554__A2 register_file\[22\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12202_ _06970_ register_file\[31\]\[6\] _06979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13182_ _07531_ _07601_ _07602_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10394_ _03830_ _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08222__A3 _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10565__A1 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12133_ _06674_ _06929_ _06934_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16195__CLK clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12306__A2 _07050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13503__A1 _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12064_ _06892_ net20 _06893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10317__A1 _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11015_ _06228_ _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_78_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12080__I _06873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15256__A1 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_92_clk_I clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15823_ _00211_ clknet_leaf_127_clk register_file\[26\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15754_ _00142_ clknet_leaf_95_clk register_file\[13\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11817__A1 _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12966_ _07458_ register_file\[17\]\[1\] _07460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14705_ register_file\[3\]\[12\] _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11917_ _06698_ _06799_ _06804_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12490__A1 _06999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15685_ _00073_ clknet_leaf_72_clk register_file\[28\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11293__A2 _06408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12897_ _07414_ register_file\[18\]\[5\] _07419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11424__I _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14636_ _02144_ _01811_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11848_ _06710_ _06758_ _06762_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_150_clk_I clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14231__A2 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11045__A2 _06250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14567_ _01741_ register_file\[17\]\[11\] _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11779_ _06721_ _06722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14782__A3 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16306_ _00694_ clknet_leaf_158_clk register_file\[21\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08997__A1 _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12793__A2 register_file\[20\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_clk_I clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13518_ _01038_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_179_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14498_ _02007_ _01757_ _02008_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16237_ _00625_ clknet_leaf_139_clk register_file\[23\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12255__I _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13449_ _07756_ register_file\[9\]\[22\] _07762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_165_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08749__A1 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12545__A2 register_file\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16168_ _00556_ clknet_leaf_92_clk register_file\[25\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15119_ register_file\[4\]\[17\] _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ _04307_ _04310_ _03817_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16099_ _00487_ clknet_leaf_14_clk register_file\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15495__A1 _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07972__A2 _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07941_ _03274_ register_file\[14\]\[25\] _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10308__A1 _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09174__A1 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07872_ _03206_ _02958_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15247__A1 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08921__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09611_ _04855_ register_file\[19\]\[15\] _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_103_clk_I clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09542_ _03810_ _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11808__A1 _06670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12481__A1 _07150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09473_ _04582_ register_file\[24\]\[13\] _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_90_clk clknet_5_14__leaf_clk clknet_leaf_90_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_149_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11334__I _06155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08424_ _03751_ _03657_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09229__A2 register_file\[17\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14222__A2 register_file\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11036__A2 _06243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15250__B _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16068__CLK clknet_leaf_313_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08355_ register_file\[7\]\[31\] _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12233__A1 _06995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08988__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13981__A1 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08286_ _01043_ register_file\[18\]\[30\] _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10795__A1 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12536__A2 register_file\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09401__A2 register_file\[19\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_30__f_clk clknet_3_7_0_clk clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15905__CLK clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15486__A1 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14289__A2 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07963__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09165__A1 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08912__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09809_ _05117_ register_file\[22\]\[18\] _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12820_ _07250_ _07370_ _07372_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14461__A2 register_file\[24\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12751_ _07326_ register_file\[20\]\[11\] _07331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12472__A1 _07150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_81_clk clknet_5_11__leaf_clk clknet_leaf_81_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08140__A2 register_file\[26\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11702_ _06072_ _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15470_ _02968_ _02969_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12682_ _07279_ register_file\[21\]\[20\] _07285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14213__A2 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14421_ _01932_ register_file\[8\]\[9\] _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11633_ _06414_ _06616_ _06621_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08979__A1 _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12775__A2 register_file\[20\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14352_ _01603_ register_file\[14\]\[8\] _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08553__I _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11564_ _06579_ register_file\[11\]\[23\] _06580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13303_ _07631_ register_file\[14\]\[28\] _07674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12075__I _06862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10515_ _05750_ register_file\[10\]\[28\] _05814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14283_ register_file\[3\]\[7\] _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11495_ _06495_ register_file\[12\]\[28\] _06538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12527__A2 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16022_ _00410_ clknet_leaf_237_clk register_file\[6\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13234_ _07630_ _07633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10446_ _05728_ _05745_ _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10377_ _05609_ register_file\[31\]\[26\] _05678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13165_ _07590_ register_file\[15\]\[4\] _07592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12803__I _07361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12116_ _06658_ _06922_ _06924_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13096_ _07519_ _07544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12047_ _06878_ net13 _06883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08903__A1 _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10710__A1 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15806_ _00194_ clknet_leaf_28_clk register_file\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13998_ _01249_ register_file\[10\]\[4\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15737_ _00125_ clknet_leaf_262_clk register_file\[27\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11266__A2 _06384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12949_ _07443_ register_file\[18\]\[27\] _07449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11154__I _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_72_clk clknet_5_10__leaf_clk clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15668_ _00056_ clknet_leaf_210_clk register_file\[2\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11018__A2 register_file\[28\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14619_ _02121_ _02128_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14465__I _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15599_ _03087_ _03096_ _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08140_ _03229_ register_file\[26\]\[28\] _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12766__A2 _07336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16360__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08071_ _03320_ register_file\[23\]\[27\] _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12518__A2 _07174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13715__A1 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13191__A2 _07601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12713__I _06159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15468__A1 _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08973_ _04293_ _04294_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09147__A1 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14140__A1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07924_ _03256_ _03009_ _03257_ _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07855_ _03186_ _03189_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10701__A1 _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13544__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07786_ _03119_ _03121_ _02953_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ _04633_ register_file\[1\]\[13\] _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12454__A1 _07138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_63_clk clknet_5_9__leaf_clk clknet_leaf_63_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08122__A2 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09456_ _04630_ register_file\[2\]\[12\] _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12206__A1 _06980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11009__A2 _06229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08407_ _03706_ register_file\[26\]\[31\] _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_71_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07881__A1 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09387_ _04630_ register_file\[2\]\[11\] _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12757__A2 _07329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13954__A1 _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08338_ _00995_ _03666_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08373__I _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09622__A2 register_file\[9\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10768__A1 _06042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08425__A3 _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08269_ _03598_ _01052_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10300_ _05600_ _05601_ _05602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12509__A2 _07167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11280_ _06085_ _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14324__B _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10231_ _05532_ _05533_ _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13182__A2 _07601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11193__A1 _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08322__B _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output79_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10162_ _05397_ register_file\[8\]\[23\] _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10940__A1 _06189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11239__I _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14131__A1 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10143__I _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14970_ _02474_ register_file\[24\]\[16\] _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10093_ _05397_ register_file\[28\]\[22\] _05398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13921_ _01437_ _01258_ _01438_ _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12693__A1 _07290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11496__A2 _06534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08361__A2 _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13852_ _01370_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12803_ _07361_ _07362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12445__A1 _07087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16571_ _00959_ clknet_leaf_285_clk register_file\[29\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11248__A2 _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13783_ _01216_ register_file\[23\]\[2\] _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_54_clk clknet_5_8__leaf_clk clknet_leaf_54_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10995_ _06221_ register_file\[28\]\[2\] _06224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09310__A1 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15522_ _02934_ register_file\[11\]\[22\] _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12996__A2 register_file\[17\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12734_ _07244_ _07312_ _07320_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16383__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15453_ _01092_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12665_ _07267_ register_file\[21\]\[15\] _07273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11702__I _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14404_ _01915_ _01832_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11616_ _06398_ _06609_ _06611_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15384_ _02876_ _02884_ _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12596_ _07026_ _07222_ _07224_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08416__A3 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14335_ _01838_ _01847_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11547_ _06565_ register_file\[11\]\[16\] _06570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11420__A2 _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14266_ _01605_ register_file\[15\]\[7\] _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11478_ _06419_ _06527_ _06528_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16005_ _00393_ clknet_leaf_313_clk register_file\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13217_ _07619_ register_file\[15\]\[25\] _07623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10429_ _03799_ _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14197_ _01711_ _01538_ _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11184__A1 _06078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13148_ _06162_ _07580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10931__A1 _06069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14122__A1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13079_ _07519_ _07532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14673__A2 register_file\[8\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10988__I _06218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11487__A2 _06527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13364__I _07689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08352__A2 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09063__B _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14425__A2 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12436__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09301__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09310_ _04494_ register_file\[11\]\[10\] _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12987__A2 _07466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10998__A1 _06225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09241_ _04558_ register_file\[28\]\[9\] _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15750__CLK clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11612__I _06601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12739__A2 register_file\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09172_ _04489_ _04490_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08123_ _03380_ register_file\[2\]\[27\] _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11411__A2 register_file\[26\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16106__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08054_ _03386_ _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13164__A2 _07584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12911__A2 register_file\[18\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10922__A1 _06050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16256__CLK clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07981__B _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _04276_ _04277_ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input30_I new_value[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07907_ _03237_ _03240_ _03075_ _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12675__A1 _07279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11478__A2 _06527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10898__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08887_ _04202_ _04209_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08343__A2 _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07838_ _03171_ _03089_ _03172_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10150__A2 register_file\[31\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_36_clk clknet_5_6__leaf_clk clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09508_ _04689_ register_file\[30\]\[13\] _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12978__A2 _07466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10780_ _06064_ _06052_ _06066_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09843__A2 register_file\[31\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09439_ _03765_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12618__I _06036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11650__A2 _06630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12450_ _07134_ _07137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_36_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11401_ _06476_ register_file\[26\]\[22\] _06482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11402__A2 _06479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12381_ _07094_ register_file\[24\]\[4\] _07096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14120_ _00994_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_153_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11332_ _06368_ register_file\[19\]\[28\] _06439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14352__A1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14051_ _01478_ register_file\[30\]\[5\] _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11263_ _06063_ _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11166__A1 _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08052__B _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13002_ _07271_ _07480_ _07481_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12902__A2 _07418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10214_ _05515_ _05516_ _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11194_ _06095_ _06344_ _06345_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10913__A1 _06037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10145_ _03823_ _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15623__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10076_ _05114_ register_file\[16\]\[22\] _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14953_ _02456_ _02458_ _02127_ _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12666__A1 _07271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09531__A1 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13904_ _01420_ _01421_ _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14884_ _01058_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12418__A1 _07116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13835_ _00998_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_clk clknet_5_3__leaf_clk clknet_leaf_27_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16554_ _00942_ clknet_leaf_105_clk register_file\[29\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12969__A2 _07456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13091__A1 _07538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13766_ _01276_ _01285_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10978_ _06156_ _06206_ _06211_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15505_ _03003_ register_file\[28\]\[22\] _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07845__A1 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12717_ _07232_ register_file\[21\]\[31\] _07309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16485_ _00873_ clknet_leaf_61_clk register_file\[15\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12528__I _07182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13697_ _01216_ register_file\[23\]\[1\] _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16129__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15436_ _01138_ _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12648_ _07255_ register_file\[21\]\[10\] _07261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09598__A1 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15367_ _02867_ _02620_ _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12579_ _07009_ _07208_ _07214_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09837__I _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14318_ _01830_ _01488_ _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08270__A1 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15298_ _02798_ _02799_ _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13359__I _07678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16279__CLK clknet_leaf_197_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13146__A2 register_file\[16\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14249_ _01739_ _01762_ _01506_ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11157__A1 _06021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09770__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08810_ _04061_ register_file\[28\]\[3\] _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _05098_ _05099_ _05100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14646__A2 _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10380__A2 _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08741_ _04064_ _04065_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11607__I _06593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09522__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08672_ _03905_ register_file\[10\]\[1\] _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12409__A1 _07109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11880__A2 register_file\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_18_clk clknet_5_2__leaf_clk clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08089__A1 _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09521__B _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07820__I _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07836__A1 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11632__A2 register_file\[10\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09224_ _04540_ _04541_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13978__B _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09589__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14582__A1 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09155_ _04473_ register_file\[8\]\[8\] _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08106_ _03435_ _03436_ _03437_ _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09086_ _04404_ _04405_ _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13137__A2 register_file\[16\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08037_ _03366_ _03368_ _03369_ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_163_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14885__A2 register_file\[25\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15646__CLK clknet_leaf_304_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08013__A1 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09761__A1 _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09988_ _05287_ _05294_ _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14637__A2 register_file\[27\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12648__A1 _07255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08939_ _04258_ _04260_ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15796__CLK clknet_leaf_172_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09513__A1 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08316__A2 register_file\[9\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11950_ _06652_ _06816_ _06824_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11320__A1 _06429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10123__A2 register_file\[14\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10901_ _06026_ register_file\[30\]\[31\] _06165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11881_ _06662_ _06778_ _06783_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13620_ _01093_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10832_ _06025_ _06109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13073__A1 _07527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09816__A2 register_file\[6\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13551_ _01071_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11623__A2 _06609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12820__A1 _07250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10763_ _06042_ register_file\[30\]\[5\] _06053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11252__I _06049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12502_ _07011_ _07167_ _07168_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16270_ _00658_ clknet_leaf_153_clk register_file\[22\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13482_ net7 net8 _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10694_ _03841_ register_file\[5\]\[31\] _05990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15221_ _02474_ register_file\[16\]\[19\] _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12433_ _07123_ register_file\[24\]\[25\] _07127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07886__B _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16421__CLK clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11387__A1 _06469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15152_ _02321_ register_file\[22\]\[18\] _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12364_ _07034_ _07042_ _07084_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08252__A1 _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14103_ _01618_ _01271_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13128__A2 _07556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11315_ _06367_ _06427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15083_ _02586_ register_file\[20\]\[17\] _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12295_ _06965_ _07040_ _07044_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11139__A1 _06148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14034_ _00999_ _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08004__A1 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11246_ _06370_ _06378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12887__A1 _07237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09752__A1 _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11177_ _06064_ _06330_ _06335_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10362__A2 register_file\[5\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10128_ _05228_ register_file\[9\]\[22\] _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15985_ _00373_ clknet_leaf_229_clk register_file\[7\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11427__I _06497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08307__A2 register_file\[29\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13300__A2 _07670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10059_ _05355_ _05364_ _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14936_ _01161_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10114__A2 register_file\[7\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14867_ register_file\[5\]\[14\] _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13818_ _01336_ _01117_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13064__A1 _07518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08736__I _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14798_ _02297_ _02305_ _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10487__B _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16537_ _00925_ clknet_leaf_241_clk register_file\[14\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11614__A2 _06609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12258__I _06129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13749_ _01162_ _01268_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12811__A1 _07366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11162__I _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16468_ _00856_ clknet_leaf_167_clk register_file\[16\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13367__A2 register_file\[29\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15419_ _02673_ register_file\[29\]\[21\] _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16399_ _00787_ clknet_leaf_144_clk register_file\[18\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11378__A1 _06400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15669__CLK clknet_leaf_224_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08243__A1 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10050__A1 _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13089__I _07506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14316__A1 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_7_clk clknet_5_1__leaf_clk clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09911_ _05215_ _05218_ _04675_ _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12878__A1 _07308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09743__A1 _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09842_ _05082_ register_file\[30\]\[18\] _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12721__I _07311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11550__A1 _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07815__I _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09773_ _05082_ register_file\[6\]\[17\] _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11337__I _06159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15292__A2 _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08724_ _03861_ register_file\[5\]\[2\] _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11302__A1 _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08655_ _03979_ _03980_ _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15044__A2 register_file\[2\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13055__A1 _07514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08586_ _03912_ _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10397__B _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11072__I _06270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08482__A1 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15479__I _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09207_ _04523_ _04524_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13358__A2 _07704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11369__A1 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09138_ _04455_ _04456_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08234__A1 _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16594__CLK clknet_leaf_176_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12030__A2 _06864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14307__A1 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10041__A1 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09982__A1 _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__A2 register_file\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09069_ _04386_ _04388_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10592__A2 register_file\[7\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11100_ _06283_ register_file\[27\]\[11\] _06288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12080_ _06873_ _06902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_46_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12869__A1 _07395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13727__I _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11031_ _06100_ _06243_ _06245_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11541__A1 _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output61_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15770_ _00158_ clknet_leaf_255_clk register_file\[13\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12982_ _07252_ _07466_ _07469_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13294__A1 _07667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14721_ _02227_ _02228_ _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11933_ _06767_ register_file\[6\]\[31\] _06813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11844__A2 _06758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14652_ _02158_ _02160_ _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11864_ _06770_ register_file\[6\]\[2\] _06773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13046__A1 _07502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08556__I _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13603_ _01123_ register_file\[10\]\[0\] _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10815_ _06094_ _06095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14794__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13597__A2 _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14583_ _02084_ _02092_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11795_ _06726_ register_file\[7\]\[6\] _06732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16322_ _00710_ clknet_leaf_60_clk register_file\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13534_ _00993_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_186_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10746_ _06037_ _06027_ _06038_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15811__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15389__I _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10280__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13349__A2 _07697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14546__A1 _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16253_ _00641_ clknet_leaf_34_clk register_file\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13465_ _07727_ register_file\[9\]\[29\] _07771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10677_ _05965_ _05972_ _05973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15204_ _02371_ _02706_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12416_ _07116_ register_file\[24\]\[18\] _07117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08225__A1 _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16184_ _00572_ clknet_leaf_191_clk register_file\[25\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12021__A2 _06864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13396_ _07730_ register_file\[9\]\[0\] _07731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09973__A1 _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15135_ _02629_ _02638_ _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08776__A2 register_file\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12347_ _07038_ _07075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15961__CLK clknet_leaf_257_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14849__A2 register_file\[10\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11780__A1 _06722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15066_ _02321_ register_file\[30\]\[17\] _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12278_ _06155_ _07032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_190_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13637__I _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14017_ register_file\[5\]\[4\] _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11229_ _06319_ register_file\[13\]\[31\] _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16317__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15274__A2 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13285__A1 _07660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12088__A2 _06902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15968_ _00356_ clknet_5_0__leaf_clk register_file\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10099__A1 _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_4_clk_I clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14919_ _02176_ register_file\[23\]\[15\] _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15899_ _00287_ clknet_leaf_265_clk register_file\[11\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16467__CLK clknet_leaf_167_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15026__A2 _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08440_ _03766_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_91_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08466__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13037__A1 _07455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13588__A2 register_file\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08371_ _03698_ _01197_ _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12260__A2 register_file\[31\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10271__A1 _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12716__I _06163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08216__A1 _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12012__A2 _06818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10023__A1 _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09964__A1 _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08767__A2 register_file\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11771__A1 _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10574__A2 register_file\[24\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13547__I _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12451__I _07137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09246__B _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07990__A3 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11523__A1 _06550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09825_ _04998_ register_file\[15\]\[18\] _05134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09756_ _04996_ register_file\[18\]\[17\] _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13276__A1 _07546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12079__A2 _06895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08707_ _04031_ register_file\[8\]\[2\] _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09687_ _04319_ _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _03798_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13028__A1 _07298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15834__CLK clknet_leaf_265_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08569_ _03878_ _03895_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10600_ _05892_ _05897_ _05898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08455__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11580_ _06442_ _06546_ _06588_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12251__A2 _07012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14528__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10531_ _03890_ register_file\[15\]\[28\] _05830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15984__CLK clknet_leaf_230_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13250_ _07518_ _07642_ _07643_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08207__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13200__A1 _07612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10462_ _05695_ register_file\[31\]\[27\] _05762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12003__A2 register_file\[5\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12201_ _06055_ _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09955__A1 _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13181_ _07598_ register_file\[15\]\[10\] _07602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10393_ _05693_ register_file\[22\]\[26\] _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11762__A1 _06708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12132_ _06933_ register_file\[3\]\[13\] _06934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13503__A2 _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12063_ _06862_ _06892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11014_ _06069_ _06229_ _06235_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15256__A2 register_file\[31\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_240_clk clknet_5_17__leaf_clk clknet_leaf_240_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15822_ _00210_ clknet_leaf_150_clk register_file\[26\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15753_ _00141_ clknet_leaf_100_clk register_file\[13\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12965_ _07230_ _07456_ _07459_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13192__I _07593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14704_ _02131_ register_file\[2\]\[12\] _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11916_ _06803_ register_file\[6\]\[23\] _06804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15684_ _00072_ clknet_leaf_70_clk register_file\[28\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12896_ _07417_ _07418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12490__A2 _07160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14635_ _02143_ _01976_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14767__A1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11847_ _06719_ register_file\[7\]\[28\] _06762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14566_ _01994_ register_file\[16\]\[11\] _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11778_ _06718_ _06721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_92_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10253__A1 _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16305_ _00693_ clknet_leaf_159_clk register_file\[21\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08997__A2 register_file\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13517_ _01037_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10729_ _06023_ _06024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_14497_ _01758_ register_file\[23\]\[10\] _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11440__I _06505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16236_ _00624_ clknet_leaf_137_clk register_file\[23\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15192__A1 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13448_ _07558_ _07759_ _07761_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09946__A1 _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16167_ _00555_ clknet_leaf_92_clk register_file\[25\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13379_ _07715_ register_file\[29\]\[26\] _07720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15118_ _02618_ _02621_ _02537_ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16098_ _00486_ clknet_leaf_14_clk register_file\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15495__A2 register_file\[25\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15707__CLK clknet_leaf_271_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15049_ _02552_ _02553_ _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07940_ _01161_ _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10308__A2 register_file\[15\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09174__A2 register_file\[14\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07871_ register_file\[5\]\[24\] _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09610_ _04853_ register_file\[18\]\[15\] _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15247__A2 register_file\[27\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_231_clk clknet_5_21__leaf_clk clknet_leaf_231_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13258__A1 _07646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15857__CLK clknet_leaf_171_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09541_ _04853_ register_file\[26\]\[14\] _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14198__I _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11808__A2 _06737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09472_ _04580_ register_file\[25\]\[13\] _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12481__A2 register_file\[23\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10492__A1 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08423_ register_file\[23\]\[31\] _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08354_ _01179_ register_file\[6\]\[31\] _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12233__A2 register_file\[31\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13430__A1 _07749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14147__B _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10244__A1 _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_298_clk clknet_5_4__leaf_clk clknet_leaf_298_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08988__A2 register_file\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13981__A2 register_file\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08285_ _01069_ register_file\[19\]\[30\] _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10795__A2 register_file\[30\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11992__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_272_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09937__A1 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14930__A1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11744__A1 _06687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15486__A2 register_file\[21\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_287_clk_I clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09165__A2 register_file\[27\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15238__A2 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09808_ _03827_ _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_222_clk clknet_5_21__leaf_clk clknet_leaf_222_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_210_clk_I clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13249__A1 _07638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14997__A1 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09739_ _04781_ register_file\[10\]\[17\] _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12750_ _07259_ _07329_ _07330_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11701_ _06665_ _06656_ _06666_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_225_clk_I clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12681_ _07247_ _07284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_15__f_clk_I clknet_3_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14420_ _01079_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11632_ _06620_ register_file\[10\]\[18\] _06621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13421__A1 _07742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_289_clk clknet_5_5__leaf_clk clknet_leaf_289_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14351_ _01862_ _01775_ _01863_ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08979__A2 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11563_ _06542_ _06579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13972__A2 _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11260__I _06059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13302_ _07572_ _07670_ _07673_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15174__A1 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16162__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10514_ _05811_ _05812_ _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14282_ _01713_ register_file\[2\]\[7\] _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_7_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11494_ _06436_ _06534_ _06537_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16021_ _00409_ clknet_leaf_238_clk register_file\[6\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13233_ _07631_ _07632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10445_ _05737_ _05744_ _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11735__A1 _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10538__A2 _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09665__I _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13164_ _07513_ _07584_ _07591_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10376_ _05607_ register_file\[30\]\[26\] _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13187__I _07585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12115_ _06918_ register_file\[3\]\[6\] _06924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13095_ _06093_ _07543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12046_ _02038_ _06881_ _06882_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_213_clk clknet_5_23__leaf_clk clknet_leaf_213_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08903__A2 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15805_ _00193_ clknet_leaf_279_clk register_file\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14988__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13997_ _01247_ register_file\[11\]\[4\] _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15736_ _00124_ clknet_leaf_199_clk register_file\[27\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12948_ _07298_ _07446_ _07448_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10474__A1 _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15351__B _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12879_ _06023_ _03855_ _07406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15667_ _00055_ clknet_leaf_210_clk register_file\[2\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15401__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14618_ _02123_ _02126_ _02127_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_15598_ _03092_ _03095_ _02924_ _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13412__A1 _07522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16505__CLK clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12266__I _06975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14549_ _01973_ register_file\[25\]\[11\] _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09092__A1 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11974__A1 _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15165__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08070_ _03153_ register_file\[22\]\[27\] _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15577__I _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14912__A1 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16219_ _00607_ clknet_leaf_39_clk register_file\[24\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08972_ _03928_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07923_ _03010_ register_file\[23\]\[25\] _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14140__A2 register_file\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12151__A1 _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13825__I _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_204_clk clknet_5_22__leaf_clk clknet_leaf_204_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07854_ _03187_ _03188_ _03108_ _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10701__A2 register_file\[25\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14979__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07785_ _03120_ _03037_ _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16035__CLK clknet_leaf_314_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11345__I _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09524_ _04837_ register_file\[3\]\[13\] _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08658__A1 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12454__A2 register_file\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10465__A1 _05755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09455_ _04766_ _04769_ _04220_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13560__I _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08406_ _03731_ _03733_ _01170_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__16185__CLK clknet_leaf_196_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09386_ _04698_ _04701_ _04553_ _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12206__A2 _06976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13403__A1 _07734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07881__A2 register_file\[1\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08337_ register_file\[4\]\[30\] _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10768__A2 register_file\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11965__A1 _06830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08268_ _03592_ _03597_ _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_91_clk_I clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13706__A2 _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08199_ _03529_ _01156_ _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11717__A1 _06675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08189__A3 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10230_ _05397_ register_file\[8\]\[24\] _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11193__A2 register_file\[13\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12390__A1 _06980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10161_ _05395_ register_file\[9\]\[23\] _05465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10940__A2 register_file\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14131__A2 register_file\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10092_ _03802_ _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12142__A1 _06684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13920_ _01143_ register_file\[15\]\[3\] _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12693__A2 _07284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13851_ _01187_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12802_ _07358_ _07361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_90_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_164_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08649__A1 _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16570_ _00958_ clknet_leaf_253_clk register_file\[29\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13782_ _01043_ register_file\[22\]\[2\] _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12445__A2 register_file\[24\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10994_ _06033_ _06219_ _06223_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16528__CLK clknet_leaf_173_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15521_ _03019_ _02687_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12733_ _07318_ register_file\[20\]\[4\] _07320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_44_clk_I clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15452_ _02951_ _02620_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12664_ _07247_ _07272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__15395__A1 _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14403_ _01913_ _01914_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_179_clk_I clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11615_ _06606_ register_file\[10\]\[11\] _06611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09074__A1 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15383_ _02883_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12595_ _07219_ register_file\[22\]\[26\] _07224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11956__A1 _06658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14334_ _01843_ _01846_ _01671_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_59_clk_I clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11546_ _06407_ _06568_ _06569_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14265_ _01603_ register_file\[14\]\[7\] _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11477_ _06524_ register_file\[12\]\[20\] _06528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11708__A1 _06670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09395__I _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16004_ _00392_ clknet_leaf_314_clk register_file\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13216_ _07593_ _07622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10428_ _05720_ _05727_ _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14196_ _01703_ _01710_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11184__A2 _06337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12381__A1 _07094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13147_ _07578_ _07507_ _07579_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07927__A3 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10359_ _05658_ _05659_ _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10931__A2 _06178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_117_clk_I clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14122__A2 register_file\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13078_ _06071_ _07531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16058__CLK clknet_leaf_248_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12133__A1 _06674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13645__I _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12029_ _06870_ net37 _06872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13881__A1 _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10695__A1 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08352__A3 _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12436__A2 _07126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10447__A1 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15719_ _00107_ clknet_leaf_88_clk register_file\[27\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07799__B _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10998__A2 register_file\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09240_ _03900_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15386__A1 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07863__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09171_ _04213_ register_file\[12\]\[8\] _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11947__A1 _06822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08122_ _03453_ _03210_ _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15138__A1 _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08812__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08053_ _03384_ _03385_ _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07818__I _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12372__A1 _07090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10922__A2 _06178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15310__A1 _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08955_ _03988_ register_file\[27\]\[5\] _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13555__I _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07906_ _03238_ _03155_ _03239_ _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09254__B _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08886_ _04205_ _04208_ _03992_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12675__A2 register_file\[21\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input23_I new_value[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10686__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07837_ _03090_ register_file\[29\]\[24\] _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14416__A3 _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09507_ _04819_ _04820_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10438__A1 _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09438_ _04747_ _04752_ _04118_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15377__A1 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09056__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09369_ _04681_ _04684_ _04045_ _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11400_ _06422_ _06479_ _06481_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15129__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12380_ _06969_ _07088_ _07095_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11331_ _06151_ _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10610__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output91_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14050_ _01563_ _01475_ _01565_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14352__A2 register_file\[14\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11262_ _06388_ _06384_ _06389_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13001_ _07477_ register_file\[17\]\[15\] _07481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12363__A1 _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11166__A2 _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16200__CLK clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10213_ _05449_ register_file\[16\]\[24\] _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11193_ _06341_ register_file\[13\]\[15\] _06345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10913__A2 _06168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10144_ _05447_ register_file\[29\]\[23\] _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15166__B _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12115__A1 _06918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10075_ _05112_ register_file\[17\]\[22\] _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08559__I _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14952_ _02457_ _02125_ _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12666__A2 _07272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16350__CLK clknet_leaf_303_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13903_ _01242_ register_file\[9\]\[3\] _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14883_ _02057_ register_file\[24\]\[15\] _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_5_30__f_clk_I clknet_3_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15918__CLK clknet_leaf_187_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13834_ register_file\[7\]\[2\] _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12418__A2 register_file\[24\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13615__A1 _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16553_ _00941_ clknet_5_15__leaf_clk register_file\[29\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13765_ _01284_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09295__A1 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10977_ _06167_ register_file\[2\]\[29\] _06211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08098__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13091__A2 _07532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11713__I _06642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15504_ _01318_ _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12716_ _06163_ _07308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16484_ _00872_ clknet_leaf_57_clk register_file\[15\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13696_ _01047_ _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_189_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12647_ _07247_ _07260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15435_ _02934_ register_file\[11\]\[21\] _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13918__A2 _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14040__A1 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11929__A1 _06767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09598__A2 register_file\[24\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15366_ register_file\[7\]\[20\] _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12578_ _07212_ register_file\[22\]\[19\] _07214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10601__A1 _05885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12544__I _07193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14317_ _01828_ _01829_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11529_ _06390_ _06554_ _06559_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15297_ _02634_ register_file\[1\]\[19\] _02635_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14248_ _01750_ _01761_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14343__A2 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12354__A1 _07023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11157__A2 _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14179_ _01693_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08740_ _03988_ register_file\[27\]\[2\] _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08469__I _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09522__A2 register_file\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08671_ _03995_ _03996_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09802__B _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12409__A2 register_file\[24\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09286__A1 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08089__A2 register_file\[31\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11093__A1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15359__A1 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07836__A2 register_file\[28\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09223_ _04473_ register_file\[8\]\[9\] _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09589__A2 register_file\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09154_ _04124_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12593__A1 _07219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08105_ _01048_ register_file\[13\]\[27\] _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16223__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09085_ _04125_ register_file\[8\]\[7\] _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08261__A2 _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08036_ _01092_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15531__A1 _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12345__A1 _07068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11148__A2 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08013__A2 register_file\[9\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09761__A2 register_file\[20\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09987_ _05290_ _05293_ _05028_ _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08938_ _04259_ register_file\[23\]\[5\] _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12648__A2 register_file\[21\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13845__A1 _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ _04187_ _04190_ _04191_ _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11320__A2 _06420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10900_ _06163_ _06164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11880_ _06782_ register_file\[6\]\[8\] _06783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10831_ _06107_ _06108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12629__I _07234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09277__A1 _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13073__A2 register_file\[16\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14270__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13550_ _01017_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10762_ _06051_ _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_164_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12820__A2 _07370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12501_ _07164_ register_file\[23\]\[20\] _07168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13481_ _00996_ _01001_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10693_ _05973_ _05988_ _05989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15220_ _02681_ _02722_ _02473_ net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12432_ _07097_ _07126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_138_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12584__A1 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15151_ _02652_ _02318_ _02653_ _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12363_ _07039_ register_file\[25\]\[30\] _07084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14102_ register_file\[5\]\[5\] _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11314_ _06129_ _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15082_ _01318_ _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15522__A1 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12294_ _07042_ register_file\[25\]\[1\] _07044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12336__A1 _07068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11139__A2 _06307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14033_ _01202_ register_file\[24\]\[5\] _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11245_ _06040_ _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09201__A1 _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08004__A2 register_file\[30\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12887__A2 _07408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09752__A2 register_file\[17\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11176_ _06334_ register_file\[13\]\[8\] _06335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10127_ _05422_ _05431_ _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15740__CLK clknet_leaf_283_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15984_ _00372_ clknet_leaf_230_clk register_file\[7\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10058_ _05358_ _05363_ _04486_ _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14935_ _02439_ _02192_ _02440_ _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14866_ _02371_ _02372_ _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15890__CLK clknet_leaf_171_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13817_ _01335_ _01115_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09268__A1 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14797_ _02304_ _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13064__A2 _07520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11075__A1 _06271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16536_ _00924_ clknet_leaf_241_clk register_file\[14\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13748_ register_file\[4\]\[1\] _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10822__A1 _06087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16467_ _00855_ clknet_leaf_167_clk register_file\[16\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13679_ _01199_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15418_ _02586_ register_file\[28\]\[21\] _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08752__I _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16398_ _00786_ clknet_leaf_144_clk register_file\[18\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11378__A2 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09440__A1 _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15349_ _02518_ register_file\[11\]\[20\] _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08243__A2 register_file\[9\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16396__CLK clknet_leaf_140_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10050__A2 register_file\[25\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14316__A2 register_file\[17\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12327__A1 _06997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09910_ _05216_ _05217_ _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12878__A2 _07362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09841_ _05147_ _05149_ _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09743__A2 register_file\[25\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11550__A2 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09772_ _03847_ _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_154_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08723_ _04028_ _04047_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11302__A2 register_file\[19\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08654_ _03871_ register_file\[15\]\[1\] _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12449__I _07135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08585_ _03911_ _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13055__A2 register_file\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11066__A1 _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07809__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14664__I _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14004__A1 _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09206_ _04387_ register_file\[4\]\[9\] _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08662__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12566__A1 _07205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11369__A2 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09137_ _04387_ register_file\[4\]\[8\] _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09431__A1 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10041__A2 _05346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14307__A2 register_file\[29\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09068_ _04387_ register_file\[16\]\[7\] _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12318__A1 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07993__A1 _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14858__A3 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08019_ _01138_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15763__CLK clknet_leaf_177_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_13__f_clk clknet_3_3_0_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12869__A2 register_file\[1\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11030_ _06240_ register_file\[28\]\[16\] _06245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11541__A2 _06561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output54_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15283__A3 _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12981_ _07462_ register_file\[17\]\[7\] _07469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13294__A2 register_file\[14\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14720_ _01065_ _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11932_ _06714_ _06770_ _06812_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08170__A1 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14651_ _02159_ register_file\[17\]\[12\] _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11863_ _06645_ _06768_ _06772_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16269__CLK clknet_leaf_139_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13046__A2 _07505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11263__I _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10814_ _06093_ _06094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13602_ _01122_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11057__A1 _06148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14582_ _02087_ _02090_ _02091_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11794_ _06654_ _06730_ _06731_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16321_ _00709_ clknet_leaf_67_clk register_file\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10745_ _06029_ register_file\[30\]\[2\] _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13533_ _01028_ _01053_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09670__A1 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16252_ _00640_ clknet_leaf_38_clk register_file\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13464_ _07574_ _07766_ _07770_ _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10280__A2 register_file\[18\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10676_ _05968_ _05971_ _04262_ _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12557__A1 _07198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12415_ _07086_ _07116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15203_ register_file\[4\]\[18\] _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09422__A1 _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16183_ _00571_ clknet_leaf_190_clk register_file\[25\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13395_ _07729_ _07730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08225__A2 register_file\[25\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12346_ _07016_ _07071_ _07074_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15134_ _02637_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12309__A1 _07046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07984__A1 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15065_ _02567_ _02318_ _02568_ _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12277_ _07030_ _07024_ _07031_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14016_ _01531_ _01532_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11228_ _06160_ _06322_ _06364_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11159_ _06033_ _06320_ _06324_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13809__A1 _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14749__I _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15967_ _00355_ clknet_leaf_1_clk register_file\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13285__A2 register_file\[14\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10099__A2 register_file\[21\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14918_ _02173_ register_file\[22\]\[15\] _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11296__A1 _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15898_ _00286_ clknet_leaf_265_clk register_file\[11\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08161__A1 _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12269__I _06143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14849_ _02103_ register_file\[10\]\[14\] _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14234__A1 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11048__A1 _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08370_ _03692_ _03697_ _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15636__CLK clknet_leaf_210_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12796__A1 _07306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16519_ _00907_ clknet_leaf_48_clk register_file\[14\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10271__A2 register_file\[1\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14537__A2 _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12548__A1 _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08216__A2 register_file\[20\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09413__A1 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10023__A2 register_file\[5\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11220__A1 _06144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09964__A2 register_file\[24\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07975__A1 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11771__A2 _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11523__A2 register_file\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09824_ _04996_ register_file\[14\]\[18\] _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09755_ _05062_ _05064_ _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13276__A2 _07656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13563__I _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09262__B _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08706_ _03823_ _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_167_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09686_ _04996_ register_file\[6\]\[16\] _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08152__A1 _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08637_ _03955_ _03960_ _03962_ _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12179__I _06959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13028__A2 _07494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08568_ _03885_ _03892_ _03894_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14776__A2 _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16561__CLK clknet_leaf_165_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12787__A1 _07347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14394__I _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09652__A1 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08455__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08499_ _03822_ _03825_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11811__I _06721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10530_ _03887_ register_file\[14\]\[28\] _05829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12539__A1 _07190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_195_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10461_ _05693_ register_file\[30\]\[27\] _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09404__A1 _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08207__A2 register_file\[16\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12200_ _06974_ _06976_ _06977_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13180_ _07593_ _07601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09955__A2 register_file\[9\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10392_ _03778_ _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13738__I _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12131_ _06913_ _06933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11762__A2 _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12062_ _02623_ _06888_ _06891_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14700__A2 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11013_ _06233_ register_file\[28\]\[9\] _06235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12711__A1 _07232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15821_ _00209_ clknet_leaf_131_clk register_file\[26\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13473__I _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16091__CLK clknet_leaf_288_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11278__A1 _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15752_ _00140_ clknet_leaf_84_clk register_file\[13\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08567__I _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12964_ _07458_ register_file\[17\]\[0\] _07459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08143__A1 _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14703_ _02211_ _01961_ _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11915_ _06766_ _06803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15683_ _00071_ clknet_leaf_20_clk register_file\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12895_ _07409_ _07417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_166_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14634_ _02141_ _02142_ _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14767__A2 register_file\[10\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11846_ _06708_ _06758_ _06761_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12778__A1 _07288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09643__A1 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14565_ _02066_ _02074_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11777_ _06719_ _06720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_186_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16304_ _00692_ clknet_leaf_158_clk register_file\[21\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11450__A1 _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10253__A2 register_file\[24\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13516_ _00997_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10728_ _06022_ _06023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_9_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14496_ _01755_ register_file\[22\]\[10\] _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13990__A3 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16235_ _00623_ clknet_leaf_136_clk register_file\[23\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15192__A2 register_file\[13\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13447_ _07756_ register_file\[9\]\[21\] _07761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10659_ _05953_ _05954_ _05955_ _05956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_16_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11202__A1 _06348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16166_ _00554_ clknet_leaf_91_clk register_file\[25\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09946__A2 register_file\[17\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13378_ _07567_ _07718_ _07719_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12950__A1 _07300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15117_ _02619_ _02620_ _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12329_ _07061_ register_file\[25\]\[15\] _07065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16097_ _00485_ clknet_leaf_14_clk register_file\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15048_ _02217_ register_file\[1\]\[16\] _02218_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11168__I _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12702__A1 _07291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16434__CLK clknet_leaf_165_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07870_ _03203_ _03204_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13258__A2 register_file\[14\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14455__A1 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11269__A1 _06393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09540_ _03807_ _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08134__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16584__CLK clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09471_ _04780_ _04784_ _04094_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10021__B _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08422_ _03706_ register_file\[22\]\[31\] _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_149_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14758__A2 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10492__A2 register_file\[23\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12769__A1 _07278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14428__B _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08353_ _03643_ _03681_ _01200_ net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09634__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11631__I _06590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11441__A1 _06502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08284_ _03612_ _01490_ _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11992__A2 _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15183__A2 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13194__A1 _07543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09937__A2 register_file\[29\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08940__I _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14930__A2 register_file\[10\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10691__B _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13558__I _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12941__A1 _07290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11744__A2 register_file\[8\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09807_ _05113_ _05115_ _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15801__CLK clknet_leaf_261_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14389__I _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13249__A2 register_file\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10180__A1 _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07999_ _03330_ _03331_ _03168_ _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09738_ _05046_ _05047_ _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14997__A2 register_file\[20\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _04978_ _04979_ _04980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09873__A1 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15951__CLK clknet_leaf_189_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11700_ _06663_ register_file\[8\]\[9\] _06666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12680_ _06116_ _07283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11680__A1 _06649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11631_ _06590_ _06620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08428__A2 _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15013__I _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11562_ _06424_ _06575_ _06578_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14350_ _01776_ register_file\[13\]\[8\] _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11432__A1 _06498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16307__CLK clknet_leaf_209_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13301_ _07667_ register_file\[14\]\[27\] _07673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10513_ _03844_ register_file\[8\]\[28\] _05812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14281_ _01794_ _01538_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15174__A2 register_file\[31\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11493_ _06531_ register_file\[12\]\[27\] _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13185__A1 _07598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16020_ _00408_ clknet_leaf_228_clk register_file\[6\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13232_ _07630_ _07631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10444_ _05740_ _05743_ _04873_ _05744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_clk_I clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11735__A2 _06680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13163_ _07590_ register_file\[15\]\[3\] _07591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10375_ _05673_ _05675_ _05676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12114_ _06654_ _06922_ _06923_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13094_ _07541_ _07532_ _07542_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14685__A1 _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12045_ _06878_ net12 _06882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11499__A1 _06495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10171__A1 _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11716__I _06090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15804_ _00192_ clknet_leaf_276_clk register_file\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13996_ _01512_ _01427_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12999__A1 _07269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15735_ _00123_ clknet_leaf_212_clk register_file\[27\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12947_ _07443_ register_file\[18\]\[26\] _07448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09630__B _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15666_ _00054_ clknet_leaf_178_clk register_file\[2\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12878_ _07308_ _07362_ _07405_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14617_ _01169_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09616__A1 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11829_ _06748_ register_file\[7\]\[20\] _06752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08419__A2 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15597_ _03093_ _03009_ _03094_ _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13412__A2 _07738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11423__A1 _06216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14548_ _02057_ register_file\[24\]\[11\] _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09092__A2 _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14762__I _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14479_ _01650_ register_file\[31\]\[10\] _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13176__A1 _07598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16218_ _00606_ clknet_leaf_38_clk register_file\[24\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14912__A2 register_file\[18\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12923__A1 _07429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16149_ _00537_ clknet_leaf_181_clk register_file\[31\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15824__CLK clknet_leaf_169_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08971_ _04289_ _04290_ _04292_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07922_ _03007_ register_file\[22\]\[25\] _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12151__A2 register_file\[3\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07853_ _02936_ register_file\[10\]\[24\] _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10162__A1 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15974__CLK clknet_leaf_309_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07784_ register_file\[7\]\[23\] _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08107__A1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13100__A1 _07539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09523_ _03831_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09855__A1 _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09454_ _04767_ _04768_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08935__I _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10465__A2 _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11662__A1 _06444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08405_ _03732_ _01097_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09385_ _04699_ _04700_ _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_7__f_clk_I clknet_3_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13403__A2 register_file\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10217__A2 _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08336_ _03662_ _03664_ _03369_ _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11414__A1 _06436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08267_ _03594_ _03596_ _03376_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_193_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_140_clk clknet_5_26__leaf_clk clknet_leaf_140_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08198_ register_file\[3\]\[28\] _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12914__A1 _07264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11717__A2 register_file\[8\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08594__A1 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12390__A2 _07098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10160_ _05456_ _05463_ _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12920__I _07417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10091_ _05395_ register_file\[29\]\[22\] _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12142__A2 _06936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10153__A1 _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15008__I _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13850_ _01185_ _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09006__I _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12801_ _07359_ _07360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09846__A1 _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10993_ _06221_ register_file\[28\]\[1\] _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13781_ _01298_ _01036_ _01299_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13751__I _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15520_ _03018_ _02685_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11653__A1 _06627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12732_ _07241_ _07312_ _07319_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15451_ register_file\[7\]\[21\] _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12663_ _06094_ _07271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15395__A2 register_file\[19\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11271__I _06383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14402_ _01114_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11405__A1 _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11614_ _06395_ _06609_ _06610_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10208__A2 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15382_ _02881_ _02882_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09074__A2 register_file\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12594_ _07023_ _07222_ _07223_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13945__A3 _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14333_ _01844_ _01757_ _01845_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11545_ _06565_ register_file\[11\]\[15\] _06569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_131_clk clknet_5_26__leaf_clk clknet_leaf_131_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_167_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13158__A1 _07586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15847__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11476_ _06505_ _06527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14264_ _01773_ _01775_ _01777_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12905__A1 _07254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11708__A2 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16003_ _00391_ clknet_leaf_0_clk register_file\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13215_ _07565_ _07615_ _07621_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10427_ _05723_ _05726_ _04262_ _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14195_ _01705_ _01708_ _01709_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_139_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13146_ _07504_ register_file\[16\]\[30\] _07579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10358_ _05527_ register_file\[27\]\[26\] _05659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15997__CLK clknet_leaf_307_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13077_ _07529_ _07520_ _07530_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10289_ _05588_ _05590_ _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12133__A2 _06929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13330__A1 _07518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12028_ _01446_ _06864_ _06871_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10144__A1 _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13881__A2 register_file\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11892__A1 _06789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15083__A1 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_271_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13979_ _01491_ _01495_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13661__I _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15718_ _00106_ clknet_leaf_88_clk register_file\[27\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09360__B _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11644__A1 _06627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15649_ _00037_ clknet_leaf_20_clk register_file\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_286_clk_I clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13397__A1 _07502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09170_ _04211_ register_file\[13\]\[8\] _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08121_ _03447_ _03452_ _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11947__A2 register_file\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_122_clk clknet_5_24__leaf_clk clknet_leaf_122_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08812__A2 register_file\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13149__A1 _07504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08490__I _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08052_ _03051_ register_file\[1\]\[26\] _03052_ _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_175_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12372__A2 register_file\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_224_clk_I clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14649__A1 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10383__A1 _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16002__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13836__I _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15310__A2 register_file\[27\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08954_ _03986_ register_file\[26\]\[5\] _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13321__A1 _07511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07905_ _02903_ register_file\[31\]\[25\] _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10135__A1 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_189_clk clknet_5_25__leaf_clk clknet_leaf_189_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_99_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08885_ _04206_ _04207_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13872__A2 _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10260__I _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07836_ _03003_ register_file\[28\]\[24\] _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11883__A1 _06665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_239_clk_I clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10686__A2 register_file\[16\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16152__CLK clknet_leaf_190_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I new_value[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14667__I _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09828__A1 _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14821__A1 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13571__I _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13624__A2 _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09506_ _04756_ register_file\[28\]\[13\] _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11635__A1 _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08665__I _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10438__A2 register_file\[13\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09437_ _04749_ _04751_ _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15377__A2 register_file\[2\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13388__A1 _07578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09368_ _04682_ _04683_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13927__A3 _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08319_ _03647_ _01188_ _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12915__I _07409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09299_ _04416_ register_file\[24\]\[10\] _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09496__I _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11330_ _06436_ _06432_ _06437_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10610__A2 register_file\[25\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11261_ _06378_ register_file\[19\]\[7\] _06389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output84_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13000_ _07465_ _07480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10212_ _05447_ register_file\[17\]\[24\] _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12363__A2 register_file\[25\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11192_ _06329_ _06344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08031__A3 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10374__A1 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13746__I _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12650__I _06077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10143_ _03766_ _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14104__A3 _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12115__A2 register_file\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10074_ _05348_ _05379_ _05313_ net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14951_ register_file\[5\]\[15\] _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13863__A2 _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13902_ _01108_ register_file\[8\]\[3\] _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11874__A1 _06654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10677__A2 _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14882_ _02348_ _02388_ _02056_ net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13833_ _01152_ register_file\[6\]\[2\] _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09819__A1 _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14812__A1 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16552_ _00940_ clknet_leaf_85_clk register_file\[29\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11626__A1 _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13764_ _01282_ _01283_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09295__A2 register_file\[15\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10976_ _06152_ _06206_ _06210_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15503_ _02997_ _03001_ _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12715_ _07306_ _07235_ _07307_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12097__I _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16483_ _00871_ clknet_leaf_52_clk register_file\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13695_ _01043_ register_file\[22\]\[1\] _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07845__A3 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13379__A1 _07715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15434_ _01681_ _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12646_ _06072_ _07259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14040__A2 register_file\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11929__A2 register_file\[6\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104_clk clknet_5_15__leaf_clk clknet_leaf_104_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15365_ _02865_ register_file\[6\]\[20\] _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_8_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12577_ _07006_ _07208_ _07213_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14316_ _01741_ register_file\[17\]\[8\] _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11528_ _06558_ register_file\[11\]\[8\] _06559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15296_ _02462_ _02795_ _02797_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16025__CLK clknet_leaf_243_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14247_ _01754_ _01760_ _01671_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10345__I _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11459_ _06497_ _06517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12354__A2 _07078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14178_ _01092_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13656__I _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13129_ _06137_ _07567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16175__CLK clknet_leaf_144_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13303__A1 _07631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I addrS[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08670_ _03901_ register_file\[8\]\[1\] _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11865__A1 _06647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_90_clk_I clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08730__A1 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11617__A1 _06606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11093__A2 register_file\[27\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15359__A2 register_file\[15\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ _04471_ register_file\[9\]\[9\] _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09153_ _04471_ register_file\[9\]\[8\] _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12735__I _07313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12042__A1 _06878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14582__A3 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08104_ _01774_ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13790__A1 _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09084_ _04122_ register_file\[9\]\[7\] _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08035_ _03367_ _03037_ _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14334__A3 _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15531__A2 register_file\[14\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12345__A2 register_file\[25\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16518__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_clk_I clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14171__B _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09986_ _05291_ _05292_ _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14098__A2 _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08937_ _03850_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_178_clk_I clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10108__A1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13845__A2 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08868_ _04067_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_58_clk_I clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15047__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07819_ _03153_ register_file\[22\]\[24\] _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_101_clk_I clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08799_ _04122_ register_file\[25\]\[3\] _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11608__A1 _06606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10830_ _06106_ _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08395__I register_file\[31\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14270__A2 register_file\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10761_ _06028_ _06051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_73_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12500_ _07145_ _07167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_73_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10692_ _05980_ _05987_ _05988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13480_ _01000_ register_file\[17\]\[0\] _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16048__CLK clknet_leaf_230_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12431_ _07021_ _07119_ _07125_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12033__A1 _06870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08788__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12584__A2 _07215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15150_ _02403_ register_file\[21\]\[18\] _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12362_ _07032_ _07078_ _07083_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10595__A1 _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14101_ _01531_ _01616_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11313_ _06424_ _06420_ _06425_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15081_ _02580_ _02584_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12293_ _06958_ _07040_ _07043_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12336__A2 register_file\[25\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14032_ _01507_ _01548_ _01201_ net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11244_ _06375_ _06369_ _06376_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09201__A2 register_file\[27\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10347__A1 _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13476__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11175_ _06321_ _06334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15286__A1 _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10126_ _05427_ _05430_ _03876_ _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08960__A1 _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15983_ _00371_ clknet_leaf_245_clk register_file\[7\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10057_ _05360_ _05362_ _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14934_ _02193_ register_file\[13\]\[15\] _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11847__A1 _06719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14865_ register_file\[4\]\[14\] _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14100__I register_file\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13816_ _01333_ _01334_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09268__A2 register_file\[22\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14796_ _02302_ _02303_ _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16535_ _00923_ clknet_leaf_226_clk register_file\[14\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13747_ _01263_ _01265_ _01266_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10959_ _06196_ register_file\[2\]\[21\] _06201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10822__A2 register_file\[30\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16466_ _00854_ clknet_leaf_166_clk register_file\[16\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13678_ _01197_ _01104_ _01198_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__15210__A1 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15417_ _02913_ _02916_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12024__A1 _06866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12629_ _07234_ _07247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_16397_ _00785_ clknet_leaf_142_clk register_file\[18\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14564__A3 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15348_ _02848_ _02687_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09440__A2 register_file\[25\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15279_ _02773_ _02780_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15513__A2 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09864__I _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12327__A2 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09840_ _05148_ register_file\[28\]\[18\] _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12290__I _07038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08951__A1 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09771_ _05079_ _05080_ _05081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13827__A2 _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ _04038_ _04046_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11838__A1 _06755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15029__A1 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08653_ _03868_ register_file\[14\]\[1\] _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15106__I _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14010__I register_file\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08584_ _03789_ _03791_ net3 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12263__A1 _07019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11066__A2 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14004__A2 register_file\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09205_ _04385_ register_file\[5\]\[9\] _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12566__A2 register_file\[22\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13763__A1 _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09136_ _04385_ register_file\[5\]\[8\] _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09431__A2 register_file\[8\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10577__A1 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09067_ _03823_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15908__CLK clknet_leaf_62_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09774__I _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12318__A2 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08018_ _03350_ register_file\[11\]\[26\] _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07993__A2 register_file\[25\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10329__A1 _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13296__I _07641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09195__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16490__CLK clknet_leaf_114_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15268__A1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09969_ _05275_ register_file\[27\]\[20\] _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13818__A2 _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11829__A1 _06748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12980_ _07250_ _07466_ _07468_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output47_I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11931_ _06767_ register_file\[6\]\[30\] _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11544__I _06553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14650_ _01307_ _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11862_ _06770_ register_file\[6\]\[1\] _06772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13601_ _01029_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12254__A1 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10813_ net17 _06093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11057__A2 _06257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14581_ _01670_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_307_clk clknet_5_1__leaf_clk clknet_leaf_307_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11793_ _06726_ register_file\[7\]\[5\] _06731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16320_ _00708_ clknet_leaf_19_clk register_file\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13532_ _01041_ _01050_ _01052_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10744_ _06036_ _06037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_185_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16251_ _00639_ clknet_leaf_269_clk register_file\[23\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12006__A1 _06708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13463_ _07727_ register_file\[9\]\[28\] _07770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10675_ _05969_ _05970_ _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15202_ _02702_ _02704_ _02537_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12414_ _07004_ _07112_ _07115_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12557__A2 register_file\[22\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16182_ _00570_ clknet_leaf_182_clk register_file\[25\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13394_ _07726_ _07729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10568__A1 _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09422__A2 register_file\[20\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15133_ _02633_ _02636_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12345_ _07068_ register_file\[25\]\[22\] _07074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15064_ _02403_ register_file\[29\]\[17\] _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12276_ _06960_ register_file\[31\]\[28\] _07031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11719__I _06094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14015_ register_file\[4\]\[4\] _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11227_ _06319_ register_file\[13\]\[30\] _06364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08933__A1 _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11158_ _06322_ register_file\[13\]\[1\] _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10740__A1 _06029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10109_ _05148_ register_file\[4\]\[22\] _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11089_ _06056_ _06279_ _06281_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15966_ _00354_ clknet_5_1__leaf_clk register_file\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14917_ _02421_ _02257_ _02422_ _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12493__A1 _07157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11296__A2 _06408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15897_ _00285_ clknet_leaf_261_clk register_file\[11\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08249__B _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14848_ _02101_ register_file\[11\]\[14\] _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14234__A2 register_file\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11048__A2 _06250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14779_ _02033_ register_file\[6\]\[13\] _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09859__I _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16518_ _00906_ clknet_leaf_48_clk register_file\[14\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12796__A2 _07314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13993__A1 _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16363__CLK clknet_leaf_140_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16449_ _00837_ clknet_leaf_54_clk register_file\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12548__A2 _07194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09413__A2 register_file\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11220__A2 _06358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14170__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09823_ _05130_ _05131_ _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09754_ _05063_ register_file\[16\]\[17\] _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08705_ _04029_ register_file\[9\]\[2\] _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12484__A1 _07157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09685_ _04316_ _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_93_clk clknet_5_14__leaf_clk clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08152__A2 register_file\[17\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08636_ _03961_ _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15422__A1 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14225__A2 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12236__A1 _06995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08567_ _03893_ _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13984__A1 _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08498_ _03824_ register_file\[20\]\[0\] _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09652__A2 register_file\[23\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15730__CLK clknet_leaf_173_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10460_ _05757_ _05759_ _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09119_ _04367_ register_file\[29\]\[8\] _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10391_ _05690_ _05691_ _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09718__B _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15489__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12130_ _06672_ _06929_ _06932_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15880__CLK clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10970__A1 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11539__I _06545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12061_ _06885_ net19 _06891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11012_ _06064_ _06229_ _06234_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15820_ _00208_ clknet_leaf_132_clk register_file\[26\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15751_ _00139_ clknet_leaf_84_clk register_file\[13\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12475__A1 _06985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11278__A2 register_file\[19\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12963_ _07457_ _07458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11274__I _06077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_84_clk clknet_5_11__leaf_clk clknet_leaf_84_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09340__A1 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14702_ _02205_ _02210_ _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11914_ _06696_ _06799_ _06802_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15682_ _00070_ clknet_leaf_19_clk register_file\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16386__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12894_ _07244_ _07408_ _07416_ _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12227__A1 _06994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14633_ _01973_ register_file\[25\]\[12\] _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11845_ _06755_ register_file\[7\]\[27\] _06761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12778__A2 _07343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13975__A1 _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14564_ _02069_ _02073_ _01825_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11776_ _06718_ _06719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16303_ _00691_ clknet_leaf_145_clk register_file\[21\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13515_ _01035_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10727_ _03777_ net43 _06022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14495_ _02004_ _01840_ _02005_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16234_ _00622_ clknet_leaf_97_clk register_file\[23\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13446_ _07555_ _07759_ _07760_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10658_ _03922_ register_file\[1\]\[30\] _05955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16165_ _00553_ clknet_leaf_80_clk register_file\[25\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11202__A2 register_file\[13\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13377_ _07715_ register_file\[29\]\[25\] _07719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10589_ _03883_ register_file\[4\]\[29\] _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15116_ _01354_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12328_ _07049_ _07064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12950__A2 _07446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16096_ _00484_ clknet_leaf_3_clk register_file\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10961__A1 _06196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14152__A1 _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15047_ _02462_ _02549_ _02551_ _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12259_ _06959_ _07019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10713__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13664__I _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14455__A2 register_file\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12466__A1 _06974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11269__A2 _06384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15949_ _00337_ clknet_leaf_117_clk register_file\[8\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_75_clk clknet_5_10__leaf_clk clknet_leaf_75_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08134__A2 register_file\[24\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09470_ _04782_ _04783_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15404__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08421_ _03744_ _03748_ _01022_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15753__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14758__A3 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12769__A2 _07336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08352_ _03661_ _03680_ _01194_ _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08283_ _03611_ _01063_ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09398__A1 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12743__I _07313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13194__A2 _07608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12941__A2 _07439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08070__A1 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10952__A1 _06196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11359__I _06449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16259__CLK clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10704__A1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09806_ _05114_ register_file\[20\]\[18\] _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07998_ _03084_ register_file\[26\]\[26\] _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14446__A2 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09737_ _04712_ register_file\[8\]\[17\] _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12457__A1 _06967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_66_clk clknet_5_10__leaf_clk clknet_leaf_66_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08125__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09668_ _04712_ register_file\[24\]\[16\] _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12209__A1 _06983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08619_ _03800_ register_file\[25\]\[1\] _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07884__A1 _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09599_ _04909_ _04910_ _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11680__A2 _06641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11630_ _06412_ _06616_ _06619_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13957__A1 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11561_ _06572_ register_file\[11\]\[22\] _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13300_ _07570_ _07670_ _07672_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10512_ _03841_ register_file\[9\]\[28\] _05811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14280_ _01788_ _01793_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11492_ _06434_ _06534_ _06536_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09389__A1 _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13185__A2 register_file\[15\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13231_ _06023_ _03875_ _07630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__12653__I _06081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10443_ _05741_ _05742_ _05743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11196__A1 _06100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14921__A3 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07939__A2 _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13162_ _07585_ _07590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10374_ _05674_ register_file\[28\]\[26\] _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10943__A1 _06091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_5_24__f_clk_I clknet_3_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12113_ _06918_ register_file\[3\]\[5\] _06923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13093_ _07539_ register_file\[16\]\[14\] _07542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15626__CLK clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14685__A2 register_file\[13\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12044_ _06873_ _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_172_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12696__A1 _07293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13484__I _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08364__A2 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08578__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10171__A2 register_file\[26\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15803_ _00191_ clknet_leaf_275_clk register_file\[19\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13995_ _01511_ _01424_ _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_57_clk clknet_5_8__leaf_clk clknet_leaf_57_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15776__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12999__A2 _07473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15734_ _00122_ clknet_leaf_212_clk register_file\[27\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09911__B _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12946_ _07295_ _07446_ _07447_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11120__A1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12828__I _07369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15665_ _00053_ clknet_leaf_173_clk register_file\[2\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12877_ _07359_ register_file\[1\]\[31\] _07405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14616_ _02124_ _02125_ _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13948__A1 _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11828_ _06729_ _06751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_18_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15596_ _03010_ register_file\[23\]\[23\] _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14547_ _00994_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11759_ _06706_ _06704_ _06707_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12620__A1 _07239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14478_ _01904_ register_file\[30\]\[10\] _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16217_ _00605_ clknet_leaf_196_clk register_file\[24\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12563__I _07185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14373__A1 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13429_ _07538_ _07745_ _07750_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16401__CLK clknet_leaf_160_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12923__A2 register_file\[18\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16148_ _00536_ clknet_leaf_151_clk register_file\[31\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08052__A1 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10934__A1 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14125__A1 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08970_ _04291_ register_file\[1\]\[5\] _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16079_ _00467_ clknet_leaf_234_clk register_file\[4\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14676__A2 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16551__CLK clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07921_ _03253_ _03089_ _03254_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13394__I _07726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07852_ _02934_ register_file\[11\]\[24\] _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10162__A2 register_file\[8\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12439__A1 _07087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 addrD[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07783_ _02865_ register_file\[6\]\[23\] _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_48_clk clknet_5_9__leaf_clk clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08107__A2 register_file\[14\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09522_ _04630_ register_file\[2\]\[13\] _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11111__A1 _06095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09855__A2 register_file\[24\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09453_ _04494_ register_file\[15\]\[12\] _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11662__A2 _06594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08404_ register_file\[25\]\[31\] _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09384_ _04494_ register_file\[19\]\[11\] _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14600__A2 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08335_ _03663_ _01167_ _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11414__A2 _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08266_ _03595_ _03374_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15156__A3 _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13569__I _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16081__CLK clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11178__A1 _06334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08197_ _03380_ register_file\[2\]\[28\] _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14903__A3 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12914__A2 _07425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15649__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10925__A1 _06174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09791__A1 _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08594__A2 register_file\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10090_ _03799_ _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12678__A1 _07279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15799__CLK clknet_leaf_214_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09543__A1 _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08346__A2 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10153__A2 register_file\[17\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11350__A1 _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_39_clk clknet_5_7__leaf_clk clknet_leaf_39_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12800_ _07358_ _07359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13780_ _01039_ register_file\[21\]\[2\] _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11102__A1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10992_ _06021_ _06219_ _06222_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09846__A2 register_file\[17\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12731_ _07318_ register_file\[20\]\[3\] _07319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07857__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12850__A1 _07388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11653__A2 register_file\[10\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15024__I _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15450_ _02865_ register_file\[6\]\[21\] _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12662_ _07269_ _07260_ _07270_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14401_ _01911_ _01912_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11613_ _06606_ register_file\[10\]\[10\] _06610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11405__A2 _06479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15381_ _02634_ register_file\[1\]\[20\] _02635_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12602__A1 _07032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16424__CLK clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_0_clk_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12593_ _07219_ register_file\[22\]\[25\] _07223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14332_ _01758_ register_file\[23\]\[8\] _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11544_ _06553_ _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08282__A1 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13479__I _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13158__A2 register_file\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12383__I _07089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09178__B _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14263_ _01776_ register_file\[13\]\[7\] _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11475_ _06417_ _06520_ _06526_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11169__A1 _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08082__B _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16002_ _00390_ clknet_leaf_0_clk register_file\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13214_ _07619_ register_file\[15\]\[24\] _07621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12905__A2 _07418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10426_ _05724_ _05725_ _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16574__CLK clknet_leaf_305_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14194_ _01169_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10916__A1 _06041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10117__B _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13145_ _06158_ _07578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10357_ _05525_ register_file\[26\]\[26\] _05658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12669__A1 _07274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13076_ _07527_ register_file\[16\]\[9\] _07530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10288_ _05589_ register_file\[20\]\[25\] _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09534__A1 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12027_ _06870_ net36 _06871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13330__A2 _07690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10144__A2 register_file\[29\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11341__A1 _06368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15083__A2 register_file\[20\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13094__A1 _07541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13978_ _01492_ _01493_ _01494_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07940__I _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12929_ _07278_ _07432_ _07437_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15717_ _00105_ clknet_leaf_69_clk register_file\[27\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07848__A1 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12841__A1 _07381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15648_ _00036_ clknet_leaf_3_clk register_file\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15386__A3 _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14594__A1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13397__A2 _07728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15579_ _03067_ _03076_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08120_ _03449_ _03451_ _03376_ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08273__A1 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13149__A2 register_file\[16\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08051_ _03294_ _03381_ _03383_ _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08025__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09773__A1 _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15941__CLK clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11580__A1 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14649__A2 register_file\[16\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08953_ _04273_ _04274_ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09525__A1 _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07904_ _03153_ register_file\[30\]\[25\] _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13321__A2 _07680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14013__I _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08884_ _03988_ register_file\[23\]\[4\] _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10135__A2 register_file\[2\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11332__A1 _06368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07835_ _03165_ _03169_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11883__A2 _06778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13852__I _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_2_clk_I clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09505_ _04754_ register_file\[29\]\[13\] _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07839__A1 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12832__A1 _07262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11635__A2 _06616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11372__I _06457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16447__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09436_ _04750_ register_file\[11\]\[12\] _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14585__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13388__A2 _07682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14683__I _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09367_ _04409_ register_file\[15\]\[11\] _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11399__A1 _06476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08318_ _03646_ _01186_ _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08264__A1 _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09298_ _04413_ register_file\[25\]\[10\] _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12060__A2 _06888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14337__A1 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08249_ _03577_ _03578_ _01025_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14888__A2 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11260_ _06059_ _06388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12899__A1 _07414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09764__A1 _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10211_ _05480_ _05514_ _05313_ net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11191_ _06091_ _06337_ _06343_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11571__A1 _06579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10374__A2 register_file\[28\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output77_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10142_ _05412_ _05446_ _05313_ net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15301__A3 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15019__I _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08319__A2 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10073_ _05365_ _05378_ _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14950_ _02371_ _02455_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11323__A1 _06427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13901_ _01397_ _01418_ _01105_ _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_14881_ _02366_ _02387_ _02054_ _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11874__A2 _06778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15065__A2 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13832_ _01341_ _01350_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13076__A1 _07527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14812__A2 register_file\[29\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16551_ _00939_ clknet_leaf_85_clk register_file\[29\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12378__I _07089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13763_ _01186_ register_file\[1\]\[1\] _01188_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11626__A2 _06616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10975_ _06167_ register_file\[2\]\[28\] _06210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15502_ _02999_ _03000_ _02751_ _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12714_ _07232_ register_file\[21\]\[30\] _07307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16482_ _00870_ clknet_leaf_53_clk register_file\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13694_ _01212_ _01036_ _01213_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15814__CLK clknet_leaf_107_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15368__A3 _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_0__f_clk clknet_3_0_0_clk clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15433_ _02932_ _02687_ _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13379__A2 register_file\[29\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12645_ _07257_ _07248_ _07258_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14576__A1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14593__I _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09687__I _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15364_ _01178_ _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08255__A1 _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12576_ _07212_ register_file\[22\]\[18\] _07213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14315_ _01572_ register_file\[16\]\[8\] _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11527_ _06545_ _06558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15295_ _02796_ _02715_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15964__CLK clknet_leaf_293_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14246_ _01756_ _01757_ _01759_ _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11458_ _06400_ _06513_ _06516_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15540__A3 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10409_ _05707_ _05708_ _05709_ _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_14177_ _01603_ register_file\[14\]\[6\] _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11389_ _06469_ register_file\[26\]\[17\] _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11562__A1 _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13128_ _07565_ _07556_ _07566_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07781__A3 _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13059_ _07516_ _07505_ _07517_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14768__I _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11865__A2 _06768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13672__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08766__I _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13067__A1 _07522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12288__I _07038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11617__A2 register_file\[10\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12814__A1 _07244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11192__I _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10310__B _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ _04522_ _04538_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14567__A1 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11920__I _06777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14031__A3 _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09152_ _03840_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12042__A2 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08103_ _03356_ register_file\[12\]\[27\] _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09083_ _04384_ _04402_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08034_ register_file\[7\]\[26\] _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13847__I register_file\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09746__A1 _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11553__A1 _06414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09985_ _05025_ register_file\[15\]\[20\] _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11367__I _06449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15295__A2 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08936_ _04257_ register_file\[22\]\[5\] _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10108__A2 register_file\[5\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08867_ _04188_ _04189_ _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07818_ _01071_ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13058__A1 _07514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08798_ _03860_ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15598__A3 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15837__CLK clknet_leaf_279_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12198__I _06975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11608__A2 register_file\[10\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12805__A1 _07230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10760_ _06049_ _06050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08485__A1 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14558__A1 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09419_ _04732_ _04733_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10691_ _05983_ _05986_ _04553_ _05987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08625__B _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12430_ _07123_ register_file\[24\]\[24\] _07125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08237__A1 _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12033__A2 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13230__A1 _07580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10044__A1 _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09985__A1 _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08788__A2 register_file\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12361_ _07039_ register_file\[25\]\[29\] _07083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13781__A2 _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14100_ register_file\[4\]\[5\] _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11312_ _06415_ register_file\[19\]\[22\] _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_270_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15080_ _02582_ _02583_ _02336_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12292_ _07042_ register_file\[25\]\[0\] _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13757__I _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09737__A1 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14031_ _01525_ _01547_ _01195_ _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11243_ _06371_ register_file\[19\]\[2\] _06376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11174_ _06060_ _06330_ _06333_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11277__I _06081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_285_clk_I clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10125_ _05428_ _05429_ _05430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_270_clk clknet_5_7__leaf_clk clknet_leaf_270_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08960__A2 register_file\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15982_ _00370_ clknet_leaf_245_clk register_file\[7\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13297__A1 _07667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10056_ _05361_ register_file\[27\]\[21\] _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14933_ _02107_ register_file\[12\]\[15\] _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11847__A2 register_file\[7\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15038__A2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13049__A1 _07509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14864_ _01530_ _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16603_ _00991_ clknet_leaf_284_clk register_file\[9\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13815_ _01242_ register_file\[9\]\[2\] _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14795_ _02217_ register_file\[1\]\[13\] _02218_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13746_ _01158_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16534_ _00922_ clknet_leaf_226_clk register_file\[14\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10958_ _06117_ _06199_ _06200_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_182_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_223_clk_I clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14549__A1 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16465_ _00853_ clknet_leaf_164_clk register_file\[16\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13677_ _01187_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10889_ _06154_ _06155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11740__I _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15210__A2 register_file\[2\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15212__I _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15416_ _02914_ _02915_ _02751_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12628_ _06049_ _07246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16396_ _00784_ clknet_leaf_140_clk register_file\[18\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12024__A2 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13221__A1 _07619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10035__A1 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15347_ _02847_ _02685_ _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12559_ _07198_ register_file\[22\]\[11\] _07203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13772__A2 _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11783__A1 _06645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_238_clk_I clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16142__CLK clknet_leaf_153_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15278_ _02776_ _02779_ _02447_ _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09728__A1 _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13667__I _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14229_ _01740_ _01742_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11535__A1 _06558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11187__I _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16292__CLK clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15277__A2 _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_261_clk clknet_5_19__leaf_clk clknet_leaf_261_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_100_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08951__A2 register_file\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09770_ _04812_ register_file\[4\]\[17\] _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_6_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13288__A1 _07558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _04041_ _04044_ _04045_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11838__A2 register_file\[7\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11915__I _06766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09900__A1 _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08652_ _03976_ _03977_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10510__A2 _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08583_ _03906_ _03909_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10040__B _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12263__A2 register_file\[31\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13460__A1 _07570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09204_ _04512_ _04521_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15201__A2 _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08219__A1 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13212__A1 _07619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12015__A2 _06214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09967__A1 _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09135_ _04445_ _04453_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14960__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13763__A2 register_file\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11774__A1 _06716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10577__A2 register_file\[27\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09066_ _04385_ register_file\[17\]\[7\] _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08017_ _01681_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11526__A1 _06388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10329__A2 register_file\[28\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09195__A2 register_file\[25\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11097__I _06278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_252_clk clknet_5_16__leaf_clk clknet_leaf_252_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09968_ _03907_ _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08919_ _04238_ _04240_ _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09899_ _04937_ register_file\[18\]\[19\] _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11829__A2 register_file\[7\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11930_ _06712_ _06806_ _06811_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14779__A1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11861_ _06638_ _06768_ _06771_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16015__CLK clknet_leaf_244_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13600_ _01120_ register_file\[11\]\[0\] _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10812_ _06091_ _06074_ _06092_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14580_ _02088_ _01757_ _02089_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12254__A2 _07012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11792_ _06729_ _06730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10265__A1 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13531_ _01051_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12656__I _06085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10743_ _06035_ _06036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15032__I _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16250_ _00638_ clknet_leaf_269_clk register_file\[23\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16165__CLK clknet_leaf_80_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13462_ _07572_ _07766_ _07769_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13203__A1 _07553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12006__A2 _06854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10674_ _03871_ register_file\[23\]\[31\] _05970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15201_ _02703_ _02620_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12413_ _07109_ register_file\[24\]\[17\] _07115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09958__A1 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16181_ _00569_ clknet_5_28__leaf_clk register_file\[25\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14871__I _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13393_ _07727_ _07728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11765__A1 _06710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10568__A2 register_file\[15\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15132_ _02634_ register_file\[1\]\[17\] _02635_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12344_ _07014_ _07071_ _07073_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_182_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13487__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12391__I _07089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15063_ _02235_ register_file\[28\]\[17\] _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12275_ _06151_ _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10904__I _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11517__A1 _06550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14014_ _01530_ _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09186__A2 _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11226_ _06156_ _06358_ _06363_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15259__A2 _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_243_clk clknet_5_17__leaf_clk clknet_leaf_243_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08933__A2 register_file\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11157_ _06021_ _06320_ _06323_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10108_ _05146_ register_file\[5\]\[22\] _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11088_ _06275_ register_file\[27\]\[6\] _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15965_ _00353_ clknet_leaf_307_clk register_file\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10039_ _05343_ _05344_ _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14916_ _02258_ register_file\[21\]\[15\] _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12493__A2 register_file\[23\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15896_ _00284_ clknet_leaf_264_clk register_file\[11\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14847_ _02353_ _02272_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_162_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13442__A1 _07756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14778_ _02278_ _02285_ _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10256__A1 _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16517_ _00905_ clknet_leaf_59_clk register_file\[14\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_42_clk_I clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13729_ _01122_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13993__A2 register_file\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15195__A1 _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16448_ _00836_ clknet_leaf_2_clk register_file\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10008__A1 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_177_clk_I clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13745__A2 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16379_ _00767_ clknet_leaf_284_clk register_file\[1\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11756__A1 _06703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_57_clk_I clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_100_clk_I clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15498__A2 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11508__A1 _06546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15682__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12181__A1 _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09822_ _05063_ register_file\[12\]\[18\] _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_234_clk clknet_5_20__leaf_clk clknet_leaf_234_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08924__A2 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_115_clk_I clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09753_ _03802_ _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16038__CLK clknet_leaf_309_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08704_ _03820_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14021__I _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09684_ _04993_ _04994_ _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12484__A2 register_file\[23\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13681__A1 _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08635_ _03912_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14956__I _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15422__A2 register_file\[31\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16188__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08566_ _03792_ net5 _03793_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12236__A2 register_file\[31\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13433__A1 _07749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12476__I _07145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13984__A2 register_file\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08497_ _03823_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15186__A1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14933__A1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13736__A2 _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09118_ _04403_ _04437_ _04298_ net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10390_ _05425_ register_file\[20\]\[26\] _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08612__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15489__A2 register_file\[23\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ _03772_ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10724__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10970__A2 _06206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12060_ _02539_ _06888_ _06890_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12172__A1 _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11011_ _06233_ register_file\[28\]\[8\] _06234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_225_clk clknet_5_21__leaf_clk clknet_leaf_225_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15110__A1 _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08391__A3 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15750_ _00138_ clknet_leaf_83_clk register_file\[13\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08679__A1 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12962_ _07454_ _07457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12475__A2 _07146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09025__I _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14701_ _02207_ _02209_ _02127_ _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11913_ _06796_ register_file\[6\]\[22\] _06802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15681_ _00069_ clknet_leaf_19_clk register_file\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12893_ _07414_ register_file\[18\]\[4\] _07416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15413__A2 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14632_ _02057_ register_file\[24\]\[12\] _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11844_ _06706_ _06758_ _06760_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12227__A2 _06988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13424__A1 _07534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14563_ _02070_ _01906_ _02072_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11775_ _06266_ _03913_ _06718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13975__A2 register_file\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11986__A1 _06844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16302_ _00690_ clknet_leaf_145_clk register_file\[21\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13514_ _01034_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10726_ _06020_ _06021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14494_ _01841_ register_file\[21\]\[10\] _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16233_ _00621_ clknet_leaf_95_clk register_file\[23\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14924__A1 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13445_ _07756_ register_file\[9\]\[20\] _07760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10657_ _03832_ register_file\[3\]\[30\] _05954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11738__A1 _06687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16164_ _00552_ clknet_leaf_75_clk register_file\[25\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13376_ _07689_ _07718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10588_ _03880_ register_file\[5\]\[29\] _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12327_ _06997_ _07057_ _07063_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15115_ register_file\[7\]\[17\] _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16095_ _00483_ clknet_leaf_3_clk register_file\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10961__A2 register_file\[2\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15046_ _02550_ _02300_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14152__A2 register_file\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12258_ _06129_ _07018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08104__I _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12163__A1 _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_216_clk clknet_5_23__leaf_clk clknet_leaf_216_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_123_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11209_ _06348_ register_file\[13\]\[22\] _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12189_ _06040_ _06969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11910__A1 _06691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10713__A2 register_file\[15\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15101__A1 _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08382__A3 _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15948_ _00336_ clknet_leaf_117_clk register_file\[8\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12466__A2 _07146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13663__A1 _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16330__CLK clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15381__B _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15879_ _00267_ clknet_leaf_109_clk register_file\[11\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13680__I _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15404__A2 register_file\[23\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14207__A3 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08420_ _03745_ _03747_ _01159_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07893__A2 _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10229__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08351_ _03672_ _03679_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11977__A1 _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15168__A1 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08282_ _03609_ _03610_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14725__B _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14915__A1 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09819__B _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09398__A2 register_file\[16\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14391__A2 _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10952__A2 register_file\[2\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14143__A2 _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14460__B _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12154__A1 _06696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_207_clk clknet_5_22__leaf_clk clknet_leaf_207_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11901__A1 _06789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09805_ _03772_ _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input39_I new_value[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07997_ _02998_ register_file\[27\]\[26\] _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09736_ _04710_ register_file\[9\]\[17\] _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12457__A2 _07136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09667_ _04710_ register_file\[25\]\[16\] _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13590__I _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08618_ _03939_ _03942_ _03943_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12209__A2 register_file\[31\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09598_ _04712_ register_file\[24\]\[15\] _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13406__A1 _07516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08549_ _03875_ _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13957__A2 register_file\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11968__A1 _06670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15159__A1 _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11560_ _06422_ _06575_ _06577_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10511_ _05794_ _05809_ _05810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14906__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11491_ _06531_ register_file\[12\]\[26\] _06536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13230_ _07580_ _07586_ _07629_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09389__A2 register_file\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10442_ _05609_ register_file\[15\]\[27\] _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14382__A2 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12393__A1 _06982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11196__A2 _06344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16203__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13161_ _07511_ _07584_ _07589_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10373_ _03900_ _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08061__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10943__A2 _06185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12112_ _06921_ _06922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15331__A1 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13092_ _06089_ _07541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12145__A1 _06686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12043_ _01955_ _06874_ _06880_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09010__A1 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12696__A2 _07284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16353__CLK clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15802_ _00190_ clknet_leaf_276_clk register_file\[19\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13994_ _01509_ _01510_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10459__A1 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15733_ _00121_ clknet_leaf_211_clk register_file\[27\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12945_ _07443_ register_file\[18\]\[25\] _07447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11120__A2 _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08808__B _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15664_ _00052_ clknet_leaf_173_clk register_file\[2\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12876_ _07306_ _07362_ _07404_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14615_ _01166_ _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09077__A1 _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11827_ _06689_ _06744_ _06750_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14070__A1 _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15595_ _03007_ register_file\[22\]\[23\] _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14546_ _02012_ _02055_ _02056_ net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11758_ _06699_ register_file\[8\]\[26\] _06707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12620__A2 _07233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10709_ _03880_ register_file\[13\]\[31\] _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14477_ _01985_ _01901_ _01987_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09639__B _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11689_ _06055_ _06658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16216_ _00604_ clknet_leaf_196_clk register_file\[24\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14373__A2 register_file\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13428_ _07749_ register_file\[9\]\[13\] _07750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12065__B _06893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16147_ _00535_ clknet_leaf_151_clk register_file\[31\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13359_ _07678_ _07708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08052__A2 register_file\[1\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10934__A2 _06185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14125__A2 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16078_ _00466_ clknet_leaf_246_clk register_file\[4\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07920_ _03090_ register_file\[21\]\[25\] _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15029_ _02450_ register_file\[6\]\[16\] _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_9_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10698__A1 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07851_ _03185_ _03104_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15720__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 addrD[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07782_ _03110_ _03117_ _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12439__A2 register_file\[24\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09521_ _04829_ _04834_ _04002_ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11111__A2 _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09452_ _04492_ register_file\[14\]\[12\] _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07866__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15870__CLK clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08403_ _03701_ register_file\[24\]\[31\] _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09383_ _04492_ register_file\[18\]\[11\] _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09068__A1 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13939__A2 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08334_ register_file\[7\]\[30\] _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_178_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14455__B _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10622__A1 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16226__CLK clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08265_ register_file\[5\]\[29\] _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08291__A2 _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15130__I _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15561__A1 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14364__A2 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08196_ _03526_ _03210_ _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11178__A2 register_file\[13\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12375__A1 _06965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10925__A2 register_file\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16376__CLK clknet_leaf_240_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12127__A1 _06926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12678__A2 register_file\[21\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09543__A2 register_file\[27\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10689__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14419__A3 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11350__A2 register_file\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15092__A3 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09719_ _05019_ _05029_ _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10991_ _06221_ register_file\[28\]\[0\] _06222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11102__A2 register_file\[27\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12730_ _07313_ _07318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07857__A2 register_file\[13\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12850__A2 register_file\[1\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12661_ _07267_ register_file\[21\]\[14\] _07270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09059__A1 _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10861__A1 _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14052__A1 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14400_ _01741_ register_file\[17\]\[9\] _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11612_ _06601_ _06609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_93_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12592_ _07193_ _07222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15380_ _02877_ _02878_ _02880_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12602__A2 _07222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_19__f_clk clknet_3_4_0_clk clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10613__A1 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12664__I _07247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14331_ _01755_ register_file\[22\]\[8\] _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11543_ _06405_ _06561_ _06567_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14262_ _01134_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11474_ _06524_ register_file\[12\]\[19\] _06526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11169__A2 register_file\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12366__A1 _07036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13213_ _07562_ _07615_ _07620_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16001_ _00389_ clknet_leaf_0_clk register_file\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10425_ _05527_ register_file\[23\]\[27\] _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14193_ _01706_ _01707_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10916__A2 _06168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13144_ _07576_ _07568_ _07577_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10356_ _05655_ _05656_ _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13709__B _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12118__A1 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15743__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09194__B _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13075_ _06067_ _07529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10287_ _03863_ _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12669__A2 _07272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13866__A1 _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12026_ _06865_ _06870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09534__A2 register_file\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15607__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15893__CLK clknet_leaf_216_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09298__A1 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13094__A2 _07532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14291__A1 _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13977_ _01075_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11743__I _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15716_ _00104_ clknet_leaf_70_clk register_file\[27\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12928_ _07436_ register_file\[18\]\[18\] _07437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A2 register_file\[9\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12841__A2 register_file\[1\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16249__CLK clknet_leaf_193_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15647_ _00035_ clknet_leaf_3_clk register_file\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12859_ _07358_ _07395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14594__A2 register_file\[10\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15578_ _03071_ _03074_ _03075_ _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10604__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14529_ register_file\[5\]\[10\] _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09369__B _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16399__CLK clknet_leaf_144_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _03382_ _03132_ _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12357__A1 _07075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09222__A1 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08025__A2 register_file\[13\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12109__A1 _06918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11580__A2 _06546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08952_ _04061_ register_file\[24\]\[5\] _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09525__A2 register_file\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07903_ _03234_ _03150_ _03236_ _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08883_ _03986_ register_file\[22\]\[4\] _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11332__A2 register_file\[19\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07834_ _03166_ _03167_ _03168_ _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09289__A1 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14282__A1 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11096__A1 _06069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09504_ _04814_ _04817_ _04057_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07839__A2 register_file\[30\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12832__A2 _07377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09435_ _03870_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09366_ _04407_ register_file\[14\]\[11\] _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14585__A2 register_file\[8\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15616__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12596__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08317_ _03644_ _03645_ _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09297_ _04610_ _04613_ _04045_ _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09279__B _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14337__A2 register_file\[8\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10071__A2 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08248_ _03352_ register_file\[10\]\[29\] _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12348__A1 _07075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14913__B _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10218__B _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15766__CLK clknet_leaf_224_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09213__A1 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08016__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08179_ _01048_ register_file\[13\]\[28\] _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12899__A2 register_file\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10210_ _05497_ _05513_ _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11020__A1 _06233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11190_ _06341_ register_file\[13\]\[14\] _06343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09764__A2 register_file\[23\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07775__A1 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11828__I _06729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10141_ _05432_ _05445_ _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10732__I _06026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10072_ _05372_ _05377_ _05378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12520__A1 _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13900_ _01408_ _01417_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09742__B _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14880_ _02379_ _02386_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13831_ _01346_ _01349_ _01148_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13076__A2 register_file\[16\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11563__I _06542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11087__A1 _06050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16550_ _00938_ clknet_leaf_85_clk register_file\[29\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13762_ _01177_ _01279_ _01281_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10974_ _06148_ _06206_ _06209_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15501_ _02667_ register_file\[26\]\[22\] _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10834__A1 _06108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12713_ _06159_ _07306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10179__I _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16481_ _00869_ clknet_leaf_22_clk register_file\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13693_ _01039_ register_file\[21\]\[1\] _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09968__I _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15432_ _02931_ _02685_ _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12644_ _07255_ register_file\[21\]\[9\] _07258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14576__A2 register_file\[21\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16541__CLK clknet_leaf_301_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12575_ _07182_ _07212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15363_ _02853_ _02863_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10907__I _06169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09452__A1 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08255__A2 register_file\[15\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14314_ _01817_ _01826_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11526_ _06388_ _06554_ _06557_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_183_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15294_ register_file\[3\]\[19\] _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12339__A1 _07009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14245_ _01758_ register_file\[23\]\[7\] _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11457_ _06510_ register_file\[12\]\[12\] _06516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11011__A1 _06233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10408_ _05640_ register_file\[1\]\[26\] _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14176_ _01689_ _01343_ _01690_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_152_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11388_ _06410_ _06472_ _06474_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11562__A2 _06575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13127_ _07563_ register_file\[16\]\[24\] _07566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10339_ _05640_ register_file\[1\]\[25\] _05641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13058_ _07514_ register_file\[16\]\[4\] _07517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12511__A1 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12009_ _06815_ register_file\[5\]\[29\] _06859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08191__A1 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13067__A2 _07520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11078__A1 _06037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12814__A2 _07360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14016__A1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09220_ _04530_ _04537_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14567__A2 register_file\[17\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12578__A1 _07212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_2_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09151_ _04454_ _04469_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15789__CLK clknet_leaf_123_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08246__A2 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08102_ _03430_ _03433_ _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15516__A1 _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09082_ _04393_ _04401_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11250__A1 _06378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08033_ _03282_ register_file\[6\]\[26\] _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_163_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09827__B _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11648__I _06601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12750__A1 _07259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11553__A2 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14024__I register_file\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09984_ _05023_ register_file\[14\]\[20\] _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08935_ _03847_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_83_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12502__A1 _07011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08866_ _03851_ register_file\[27\]\[4\] _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input21_I new_value[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08182__A1 _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07817_ _03149_ _03150_ _03151_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14255__A1 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13058__A2 register_file\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08797_ _04104_ _04120_ _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12805__A2 _07360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16564__CLK clknet_leaf_210_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14694__I _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09682__A1 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08906__B _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08692__I _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09418_ _04663_ register_file\[7\]\[12\] _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14558__A2 register_file\[29\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10690_ _05984_ _05985_ _05986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12569__A1 _07205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09349_ _04662_ _04664_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09434__A1 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__A2 register_file\[31\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13230__A2 _07586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12360_ _07030_ _07078_ _07082_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11241__A1 _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09985__A2 register_file\[15\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11311_ _06125_ _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12291_ _07041_ _07042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14030_ _01539_ _01546_ _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11242_ _06036_ _06375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09737__A2 register_file\[8\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14730__A2 _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12741__A1 _07318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11173_ _06326_ register_file\[13\]\[7\] _06333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10124_ _05361_ register_file\[15\]\[22\] _05429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15474__B _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15981_ _00369_ clknet_leaf_247_clk register_file\[7\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14494__A1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13297__A2 register_file\[14\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13773__I _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14932_ _02434_ _02437_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10055_ _03830_ _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14863_ _02367_ _02369_ _02120_ _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_5_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13049__A2 _07505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07920__A1 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16602_ _00990_ clknet_leaf_253_clk register_file\[9\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13814_ _01108_ register_file\[8\]\[2\] _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14794_ _02045_ _02298_ _02301_ _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10807__A1 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16533_ _00921_ clknet_leaf_225_clk register_file\[14\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13745_ _01264_ _01156_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10957_ _06196_ register_file\[2\]\[20\] _06200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15931__CLK clknet_leaf_265_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08816__B _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14549__A2 register_file\[25\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16464_ _00852_ clknet_leaf_166_clk register_file\[16\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11480__A1 _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13676_ _01005_ _01030_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10888_ net32 _06154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15415_ _02667_ register_file\[26\]\[21\] _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12627_ _07244_ _07233_ _07245_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16395_ _00783_ clknet_leaf_139_clk register_file\[18\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09425__A1 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14109__I register_file\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08228__A2 _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13221__A2 register_file\[15\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10035__A2 register_file\[28\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11232__A1 _06266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15346_ _02845_ _02846_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12558_ _06987_ _07201_ _07202_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12980__A1 _07250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11783__A2 _06720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12852__I _07369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11509_ _06366_ _06544_ _06547_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15277_ _02777_ _02529_ _02778_ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12489_ _07157_ register_file\[23\]\[15\] _07161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08551__B _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14228_ _01741_ register_file\[17\]\[7\] _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09728__A2 register_file\[2\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_1_clk_I clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14721__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12732__A1 _07241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16437__CLK clknet_leaf_205_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14159_ _01654_ _01673_ _01506_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08400__A2 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14485__A1 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13288__A2 _07663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11299__A1 _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ _03876_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_79_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08164__A1 _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16587__CLK clknet_leaf_115_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08651_ _03864_ register_file\[12\]\[1\] _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09900__A2 register_file\[19\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07911__A1 _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08582_ _03908_ register_file\[7\]\[0\] _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12799__A1 _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13460__A2 _07766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15403__I _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09203_ _04515_ _04520_ _04382_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13212__A2 register_file\[15\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09134_ _04448_ _04451_ _04452_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11223__A1 _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08017__I _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15559__B _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11774__A2 _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12971__A1 _07462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09065_ _03820_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08016_ _03348_ _03104_ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11526__A2 _06554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09967_ _05273_ register_file\[26\]\[20\] _05274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14476__A1 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13593__I _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08918_ _04239_ register_file\[16\]\[5\] _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09898_ _05204_ _05205_ _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14228__A1 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08849_ _03810_ _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07902__A1 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15954__CLK clknet_leaf_216_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11860_ _06770_ register_file\[6\]\[0\] _06771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10811_ _06087_ register_file\[30\]\[14\] _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11791_ _06721_ _06729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_25_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15313__I _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11462__A1 _06517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10265__A2 register_file\[30\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13530_ _01021_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10742_ net33 _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09407__A1 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13461_ _07763_ register_file\[9\]\[27\] _07769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_5_18__f_clk_I clknet_3_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10673_ _03868_ register_file\[22\]\[31\] _05969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14400__A1 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13203__A2 _07608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15200_ register_file\[7\]\[18\] _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12412_ _07002_ _07112_ _07114_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11214__A1 _06355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16180_ _00568_ clknet_leaf_162_clk register_file\[25\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15469__B _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13754__A3 _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13392_ _07726_ _07727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14373__B _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15131_ _01370_ _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11765__A2 _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12343_ _07068_ register_file\[25\]\[21\] _07073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15062_ _02562_ _02565_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12274_ _07028_ _07024_ _07029_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14703__A2 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11288__I _06383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12714__A1 _07232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14013_ _00993_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11225_ _06319_ register_file\[13\]\[29\] _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_190_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08394__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11156_ _06322_ register_file\[13\]\[0\] _06323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10107_ _05394_ _05411_ _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10920__I _06177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11087_ _06050_ _06279_ _06280_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15964_ _00352_ clknet_leaf_293_clk register_file\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08146__A1 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10038_ _05275_ register_file\[31\]\[21\] _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14915_ _02169_ register_file\[20\]\[15\] _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14219__A1 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15895_ _00283_ clknet_leaf_217_clk register_file\[11\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14846_ _02352_ _02270_ _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12847__I _07358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14777_ _02281_ _02284_ _02030_ _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11989_ _06844_ register_file\[5\]\[20\] _06848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16516_ _00904_ clknet_leaf_59_clk register_file\[14\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11453__A1 _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10256__A2 register_file\[27\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13728_ _01247_ register_file\[11\]\[1\] _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16447_ _00835_ clknet_leaf_2_clk register_file\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10367__I _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13659_ register_file\[2\]\[0\] _01179_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_31_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10008__A2 register_file\[21\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11205__A1 _06348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16378_ _00766_ clknet_leaf_255_clk register_file\[1\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11756__A2 _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12953__A1 _07407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15329_ _02829_ _02746_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15827__CLK clknet_leaf_173_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12705__A1 _07291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08385__A1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09821_ _05061_ register_file\[13\]\[18\] _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14458__A1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15977__CLK clknet_leaf_291_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09752_ _05061_ register_file\[17\]\[17\] _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08703_ _04019_ _04027_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09683_ _04729_ register_file\[4\]\[16\] _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09885__A1 _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08634_ _03957_ _03959_ _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09637__A1 _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08565_ _03888_ _03891_ _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13433__A2 register_file\[9\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11444__A1 _06386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08496_ _03771_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_284_clk_I clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_170_clk clknet_5_28__leaf_clk clknet_leaf_170_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16602__CLK clknet_leaf_253_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13197__A1 _07605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09117_ _04423_ _04436_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09048_ _04367_ register_file\[13\]\[7\] _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_299_clk_I clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11010_ _06220_ _06233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08376__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12172__A2 _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10183__A1 _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_222_clk_I clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output52_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08128__A1 _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13121__A1 _07560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12961_ _07455_ _07456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09876__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14700_ _02208_ _02125_ _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_237_clk_I clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11912_ _06694_ _06799_ _06801_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11683__A1 _06652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15680_ _00068_ clknet_leaf_16_clk register_file\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12892_ _07241_ _07408_ _07415_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14631_ _02094_ _02140_ _02056_ net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12667__I _06099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11843_ _06755_ register_file\[7\]\[26\] _06760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09628__A1 _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13424__A2 _07745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15043__I _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11435__A1 _06502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14562_ _02071_ register_file\[31\]\[11\] _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11774_ _06716_ _06643_ _06717_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08300__A1 _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16301_ _00689_ clknet_leaf_143_clk register_file\[21\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11986__A2 register_file\[5\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13513_ _01033_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10725_ _06019_ _06020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_161_clk clknet_5_31__leaf_clk clknet_leaf_161_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14493_ _01751_ register_file\[20\]\[10\] _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15177__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16282__CLK clknet_leaf_269_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13188__A1 _07605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16232_ _00620_ clknet_leaf_93_clk register_file\[23\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13444_ _07737_ _07759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14924__A2 register_file\[8\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10656_ _03780_ register_file\[2\]\[30\] _05953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11738__A2 register_file\[8\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13498__I _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12935__A1 _07436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16163_ _00551_ clknet_leaf_65_clk register_file\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13375_ _07565_ _07711_ _07717_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08603__A2 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10587_ _05877_ _05884_ _05885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15114_ _02450_ register_file\[6\]\[17\] _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_6_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12326_ _07061_ register_file\[25\]\[14\] _07063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10410__A2 _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16094_ _00482_ clknet_leaf_299_clk register_file\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14688__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15045_ register_file\[3\]\[16\] _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12257_ _07016_ _07012_ _07017_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08367__A1 _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13360__A1 _07708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11208_ _06122_ _06351_ _06353_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12188_ _06967_ _06961_ _06968_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10174__A1 _05474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11746__I _06129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11910__A2 _06799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15101__A2 register_file\[10\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11139_ _06148_ _06307_ _06310_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15947_ _00335_ clknet_leaf_115_clk register_file\[8\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14860__A1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13961__I _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10477__A2 _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15878_ _00266_ clknet_leaf_46_clk register_file\[11\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14829_ _01075_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09619__A1 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08350_ _03678_ _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10229__A2 register_file\[9\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13966__A3 _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14792__I _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08281_ _01059_ register_file\[17\]\[30\] _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_152_clk clknet_5_30__leaf_clk clknet_leaf_152_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13179__A1 _07529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14915__A2 register_file\[20\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13718__A3 _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12926__A1 _07276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14679__A1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16005__CLK clknet_leaf_313_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15340__A2 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13351__A1 _07541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12154__A2 _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10165__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09804_ _05112_ register_file\[21\]\[18\] _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07996_ _03328_ _02912_ _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13103__A1 _07539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09735_ _05012_ _05045_ _04977_ net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14967__I _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09858__A1 _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09570__B _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09666_ _04944_ _04976_ _04977_ net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08617_ _03816_ _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_27_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09597_ _04710_ register_file\[25\]\[15\] _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11391__I _06446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14603__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13406__A2 _07728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11417__A1 _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08548_ _03874_ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_165_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11968__A2 _06833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15159__A2 register_file\[25\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_143_clk clknet_5_27__leaf_clk clknet_leaf_143_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_141_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08479_ _03777_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08914__B _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10510_ _05801_ _05808_ _05809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11490_ _06431_ _06534_ _06535_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12917__A1 _07266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10441_ _05607_ register_file\[14\]\[27\] _05741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08597__A1 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12393__A2 _07098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13160_ _07586_ register_file\[15\]\[2\] _07589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10372_ _05672_ register_file\[29\]\[26\] _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12111_ _06913_ _06921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13091_ _07538_ _07532_ _07540_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_161_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13342__A1 _07531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12145__A2 _06936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12042_ _06878_ net42 _06880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10156__A1 _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09010__A2 register_file\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_41_clk_I clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15095__A1 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15801_ _00189_ clknet_leaf_261_clk register_file\[19\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_176_clk_I clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09849__A1 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13993_ _01242_ register_file\[9\]\[4\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15732_ _00120_ clknet_leaf_177_clk register_file\[27\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12944_ _07417_ _07446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10459__A2 register_file\[28\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11656__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_56_clk_I clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15663_ _00051_ clknet_leaf_146_clk register_file\[2\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12875_ _07359_ register_file\[1\]\[30\] _07404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14614_ register_file\[5\]\[11\] _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11826_ _06748_ register_file\[7\]\[19\] _06750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15594_ _03088_ _03089_ _03091_ _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15672__CLK clknet_leaf_240_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14070__A2 register_file\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14545_ _01200_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_134_clk clknet_5_26__leaf_clk clknet_leaf_134_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11757_ _06143_ _06706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10708_ _05996_ _06003_ _06004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10631__A2 _05927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14476_ _01986_ register_file\[29\]\[10\] _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_114_clk_I clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11688_ _06654_ _06656_ _06657_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16215_ _00603_ clknet_leaf_197_clk register_file\[24\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16028__CLK clknet_leaf_293_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13427_ _07729_ _07749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10639_ _05934_ _05935_ _05936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16146_ _00534_ clknet_leaf_156_clk register_file\[31\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13358_ _07548_ _07704_ _07707_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10395__A1 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12309_ _07046_ register_file\[25\]\[7\] _07053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_129_clk_I clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15322__A2 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16077_ _00465_ clknet_leaf_247_clk register_file\[4\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13289_ _07660_ register_file\[14\]\[22\] _07666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13333__A1 _07686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15028_ _02523_ _02532_ _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11476__I _06505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13884__A2 _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11895__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07850_ _03184_ _03102_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08760__A1 _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07781_ _03113_ _03116_ _02862_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14833__A1 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 addrD[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13636__A2 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09520_ _04831_ _04833_ _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11647__A1 _06429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09451_ _04764_ _04765_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08402_ _03725_ _03729_ _01101_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09382_ _04696_ _04697_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09068__A2 register_file\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14061__A2 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08333_ _01179_ register_file\[6\]\[30\] _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_177_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_125_clk clknet_5_25__leaf_clk clknet_leaf_125_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08264_ _00995_ _03593_ _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10622__A2 register_file\[31\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08195_ _03520_ _03525_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15561__A2 register_file\[25\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08579__A1 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12375__A2 _07088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10386__A1 _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12127__A2 register_file\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13324__A1 _07513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13875__A2 _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11886__A1 _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07979_ _03063_ register_file\[19\]\[26\] _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11638__A1 _06419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09718_ _05022_ _05027_ _05028_ _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15695__CLK clknet_leaf_152_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10990_ _06220_ _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_56_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09649_ _04894_ register_file\[20\]\[15\] _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13106__I _07503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12660_ _06090_ _07269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10861__A2 _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14052__A2 register_file\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11611_ _06393_ _06602_ _06608_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12591_ _07021_ _07215_ _07221_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14330_ _01839_ _01840_ _01842_ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11542_ _06565_ register_file\[11\]\[14\] _06567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11810__A1 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15001__A1 _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14261_ _01774_ _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11473_ _06414_ _06520_ _06525_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14355__A3 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16000_ _00388_ clknet_leaf_0_clk register_file\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13212_ _07619_ register_file\[15\]\[23\] _07620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12366__A2 _07042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10424_ _05525_ register_file\[22\]\[27\] _05724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14192_ _01166_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16320__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10377__A1 _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12680__I _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13143_ _07504_ register_file\[16\]\[29\] _07577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10355_ _05589_ register_file\[24\]\[26\] _05656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07793__A2 _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12118__A2 _06922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13074_ _07526_ _07520_ _07528_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10129__A1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10286_ _05587_ register_file\[21\]\[25\] _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13866__A2 register_file\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12025_ _01358_ _06864_ _06869_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16470__CLK clknet_leaf_216_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14815__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11629__A1 _06613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13976_ _01405_ register_file\[18\]\[4\] _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09298__A2 register_file\[25\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14291__A2 _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15715_ _00103_ clknet_leaf_54_clk register_file\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12927_ _07406_ _07436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15646_ _00034_ clknet_leaf_304_clk register_file\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12858_ _07288_ _07391_ _07394_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12054__A1 _06885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11809_ _06734_ register_file\[7\]\[12\] _06740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_107_clk clknet_5_14__leaf_clk clknet_leaf_107_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15577_ _01100_ _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12789_ _07347_ register_file\[20\]\[27\] _07353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15231__I _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14528_ _01954_ _02038_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11801__A1 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10604__A2 register_file\[8\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14459_ _01949_ _01970_ _01632_ _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_122_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12357__A2 register_file\[25\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09222__A2 register_file\[9\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10368__A1 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16129_ _00517_ clknet_leaf_67_clk register_file\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13306__A1 _07576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12109__A2 register_file\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08981__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08951_ _04059_ register_file\[25\]\[5\] _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07902_ _03235_ register_file\[29\]\[25\] _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11868__A1 _06649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08882_ _04203_ _04204_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15059__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07833_ _01125_ _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14806__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_25__f_clk clknet_3_6_0_clk clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14282__A2 register_file\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09503_ _04815_ _04816_ _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11096__A2 _06279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12293__A1 _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09434_ _04748_ register_file\[10\]\[12\] _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12045__A1 _06878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09365_ _04679_ _04680_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12596__A2 _07222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08316_ _03345_ register_file\[9\]\[30\] _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09296_ _04611_ _04612_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16343__CLK clknet_leaf_197_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10285__I _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08247_ _03350_ register_file\[11\]\[29\] _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12348__A2 register_file\[25\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15297__B _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08178_ _03356_ register_file\[12\]\[28\] _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09213__A2 register_file\[21\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13596__I _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11020__A2 register_file\[28\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16493__CLK clknet_leaf_125_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10140_ _05439_ _05444_ _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13848__A2 _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10071_ _05376_ _05309_ _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08724__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12520__A2 _07174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10531__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13830_ _01347_ _01258_ _01348_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_47_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14273__A2 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11087__A2 _06279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13761_ _01280_ _01182_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10973_ _06203_ register_file\[2\]\[27\] _06209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15500_ _02998_ register_file\[27\]\[22\] _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12712_ _07304_ _07296_ _07305_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10834__A2 _06096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16480_ _00868_ clknet_leaf_6_clk register_file\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13692_ _01031_ register_file\[20\]\[1\] _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15222__A1 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14025__A2 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15431_ _02928_ _02930_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12643_ _06068_ _07257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15362_ _02856_ _02861_ _02862_ _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12574_ _07004_ _07208_ _07211_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14313_ _01821_ _01824_ _01825_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11525_ _06550_ register_file\[11\]\[7\] _06557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15293_ _02548_ register_file\[2\]\[19\] _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__15710__CLK clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12339__A2 _07064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13536__A1 _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14244_ _01096_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11456_ _06398_ _06513_ _06515_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09204__A2 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10407_ _05508_ register_file\[3\]\[26\] _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11011__A2 register_file\[28\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14175_ _01344_ register_file\[13\]\[6\] _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11387_ _06469_ register_file\[26\]\[16\] _06474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08963__A1 _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13126_ _06133_ _07565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15860__CLK clknet_leaf_175_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10338_ _03776_ _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13057_ _06044_ _07516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10269_ _05303_ register_file\[2\]\[24\] _05572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08715__A1 _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12511__A2 _07167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12008_ _06710_ _06854_ _06858_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10522__A1 _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16216__CLK clknet_leaf_196_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11754__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14264__A2 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11078__A2 _06269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13959_ _01039_ register_file\[29\]\[4\] _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09140__A1 _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16366__CLK clknet_leaf_144_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12027__A1 _06870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15629_ _00017_ clknet_leaf_135_clk register_file\[30\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12578__A2 register_file\[22\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09150_ _04461_ _04468_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13775__A1 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10589__A1 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10319__B _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08101_ _03431_ _03432_ _03108_ _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09081_ _04396_ _04399_ _04400_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11250__A2 register_file\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08032_ _03355_ _03364_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14305__I _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08954__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12750__A2 _07329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09983_ _05288_ _05289_ _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08934_ _04254_ _04255_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12502__A2 _07167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08865_ _03848_ register_file\[26\]\[4\] _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10513__A1 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07816_ _02818_ register_file\[21\]\[24\] _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08796_ _04111_ _04119_ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input14_I new_value[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09131__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15204__A1 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09417_ _04661_ register_file\[6\]\[12\] _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12495__I _07134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15733__CLK clknet_leaf_211_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12569__A2 register_file\[22\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13766__A1 _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09348_ _04663_ register_file\[23\]\[11\] _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09434__A2 register_file\[10\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15507__A2 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09279_ _04592_ _04595_ _04529_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11241__A2 _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11310_ _06422_ _06420_ _06423_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07996__A2 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12290_ _07038_ _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_147_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11241_ _06373_ _06369_ _06374_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output82_I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08945__A1 _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12741__A2 register_file\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11172_ _06056_ _06330_ _06332_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10752__A1 _06041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16239__CLK clknet_leaf_153_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_0__f_clk_I clknet_3_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10123_ _05359_ register_file\[14\]\[22\] _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15980_ _00368_ clknet_leaf_249_clk register_file\[7\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14494__A2 register_file\[21\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10054_ _05359_ register_file\[26\]\[21\] _05360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14931_ _02435_ _02436_ _02276_ _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10504__A1 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09370__A1 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08173__A2 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14862_ _02368_ _02203_ _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16389__CLK clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14246__A2 _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16601_ _00989_ clknet_leaf_257_clk register_file\[9\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13813_ _01305_ _01331_ _01105_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12257__A1 _07016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14793_ _02299_ _02300_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16532_ _00920_ clknet_leaf_174_clk register_file\[14\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10807__A2 _06074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13744_ register_file\[7\]\[1\] _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10956_ _06177_ _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_16_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16463_ _00851_ clknet_leaf_148_clk register_file\[16\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12009__A1 _06815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11480__A2 _06527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13675_ _01150_ _01192_ _01195_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_189_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10887_ _06152_ _06140_ _06153_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15414_ _02581_ register_file\[27\]\[21\] _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12626_ _07242_ register_file\[21\]\[4\] _07245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16394_ _00782_ clknet_leaf_97_clk register_file\[18\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09425__A2 register_file\[23\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15345_ _02513_ register_file\[9\]\[20\] _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12557_ _07198_ register_file\[22\]\[10\] _07202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09928__B _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11508_ _06546_ register_file\[11\]\[0\] _06547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12980__A2 _07466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15276_ _02444_ register_file\[15\]\[19\] _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12488_ _07145_ _07160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10991__A1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09189__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14227_ _01307_ _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11439_ _06497_ _06505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_99_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08936__A1 _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12732__A2 _07312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14158_ _01663_ _01672_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13109_ _06111_ _07553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14089_ _01142_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14485__A2 register_file\[17\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input6_I addrS[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12496__A1 _07164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10602__B _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08279__B _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08164__A2 register_file\[23\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08650_ _03861_ register_file\[13\]\[1\] _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08581_ _03907_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15756__CLK clknet_leaf_136_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09113__A1 _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12799__A2 _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13204__I _07593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09202_ _04517_ _04519_ _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10049__B _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09133_ _03855_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09064_ _04375_ _04383_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12971__A2 register_file\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10982__A1 _06164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08015_ _03347_ _03102_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13920__A1 _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09966_ _03904_ _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_134_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14476__A2 register_file\[29\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16531__CLK clknet_leaf_174_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08917_ _03802_ _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12487__A1 _06997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09897_ _05004_ register_file\[16\]\[19\] _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_96_clk clknet_5_15__leaf_clk clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09352__A1 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08155__A2 _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08848_ _04170_ register_file\[18\]\[4\] _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14228__A2 register_file\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07902__A2 register_file\[29\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12239__A1 _06995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08779_ _04098_ _04101_ _04102_ _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09104__A1 _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10810_ _06090_ _06091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11790_ _06652_ _06720_ _06728_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10741_ _06033_ _06027_ _06034_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13739__A1 _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13460_ _07570_ _07766_ _07768_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10672_ _05966_ _05967_ _05968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09407__A2 register_file\[30\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14400__A2 register_file\[17\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12411_ _07109_ register_file\[24\]\[16\] _07114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11214__A2 register_file\[13\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12411__A1 _07109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13391_ _06316_ _03893_ _07726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_20_clk clknet_5_2__leaf_clk clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15130_ _01185_ _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12342_ _07011_ _07071_ _07072_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10973__A1 _06203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16061__CLK clknet_leaf_300_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15061_ _02563_ _02564_ _02399_ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12273_ _07019_ register_file\[31\]\[27\] _07029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15629__CLK clknet_leaf_135_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08918__A1 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14012_ _01526_ _01528_ _01266_ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12714__A2 register_file\[21\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13911__A1 _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11224_ _06152_ _06358_ _06362_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09591__A1 _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08878__I _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11155_ _06321_ _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_150_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14467__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10106_ _05403_ _05410_ _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12478__A1 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11086_ _06275_ register_file\[27\]\[5\] _06280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15963_ _00351_ clknet_leaf_285_clk register_file\[8\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09343__A1 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15779__CLK clknet_leaf_56_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10037_ _05273_ register_file\[30\]\[21\] _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14914_ _02416_ _02419_ _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15894_ _00282_ clknet_leaf_203_clk register_file\[11\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14845_ _02350_ _02351_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15504__I _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14776_ _02282_ _02112_ _02283_ _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11988_ _06825_ _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_147_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13727_ _01119_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16515_ _00903_ clknet_leaf_22_clk register_file\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10939_ _06169_ _06189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11453__A2 register_file\[12\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13024__I _07465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13658_ _01178_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_16446_ _00834_ clknet_leaf_304_clk register_file\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12609_ _07231_ _07232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12402__A1 _06992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11205__A2 register_file\[13\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16377_ _00765_ clknet_leaf_202_clk register_file\[1\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16404__CLK clknet_leaf_173_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13589_ _00997_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14942__A3 _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_clk clknet_5_3__leaf_clk clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15328_ _02827_ _02828_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12953__A2 register_file\[18\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10964__A1 _06203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12084__B _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15259_ _02753_ _02760_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13902__A1 _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10716__A1 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09582__A1 _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09820_ _05121_ _05128_ _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14458__A2 _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09751_ _03820_ _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12469__A1 _07142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_78_clk clknet_5_10__leaf_clk clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09334__A1 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08702_ _04022_ _04025_ _04026_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08137__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09682_ _04727_ register_file\[5\]\[16\] _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11141__A1 _06152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09885__A2 register_file\[27\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _03958_ register_file\[7\]\[1\] _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07896__A1 _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13969__A1 _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08564_ _03890_ register_file\[11\]\[0\] _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09412__I _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12641__A1 _07255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11444__A2 _06506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08495_ _03821_ register_file\[21\]\[0\] _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08028__I _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13869__I _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16084__CLK clknet_leaf_230_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09116_ _04430_ _04435_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10955__A1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14146__A1 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09047_ _03766_ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_108_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08376__A2 _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11380__A1 _06469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ _05253_ _05255_ _05256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_69_clk clknet_5_10__leaf_clk clknet_leaf_69_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10242__B _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09325__A1 _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08128__A2 register_file\[1\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13121__A2 _07556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12960_ _07454_ _07455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11132__A1 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output45_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11911_ _06796_ register_file\[6\]\[21\] _06801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07887__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11683__A2 _06641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12891_ _07414_ register_file\[18\]\[3\] _07415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08647__B _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14630_ _02116_ _02139_ _02054_ _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11842_ _06703_ _06758_ _06759_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_0_clk_I clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14561_ _01649_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12632__A1 _07246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11773_ _06640_ register_file\[8\]\[31\] _06717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16300_ _00688_ clknet_leaf_139_clk register_file\[21\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13512_ _01023_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08300__A2 _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10724_ net11 _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14492_ _01999_ _02002_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16231_ _00619_ clknet_leaf_90_clk register_file\[23\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14385__A1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13443_ _07553_ _07752_ _07758_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09478__B _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10655_ _05948_ _05951_ _05028_ _05952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12935__A2 register_file\[18\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16162_ _00550_ clknet_leaf_65_clk register_file\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08064__A1 _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13374_ _07715_ register_file\[29\]\[24\] _07717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16577__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10586_ _05880_ _05883_ _03837_ _05884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10946__A1 _06095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15113_ _02607_ _02616_ _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12325_ _06994_ _07057_ _07062_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07811__A1 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16093_ _00481_ clknet_leaf_299_clk register_file\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14688__A2 register_file\[15\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15044_ _02548_ register_file\[2\]\[16\] _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12256_ _07007_ register_file\[31\]\[22\] _07017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12699__A1 _07291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11207_ _06348_ register_file\[13\]\[21\] _06353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09564__A1 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12187_ _06963_ register_file\[31\]\[2\] _06968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11371__A1 _06393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11138_ _06304_ register_file\[27\]\[27\] _06310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_6__f_clk clknet_3_1_0_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10152__B _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13019__I _07454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08119__A2 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15946_ _00334_ clknet_5_13__leaf_clk register_file\[8\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11069_ _06267_ _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11123__A1 _06117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_0_clk clknet_5_0__leaf_clk clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15877_ _00265_ clknet_leaf_63_clk register_file\[11\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12871__A1 _07359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15234__I _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14828_ _02252_ register_file\[18\]\[14\] _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12623__A1 _07242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14759_ _01932_ register_file\[8\]\[13\] _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08280_ _03306_ register_file\[16\]\[30\] _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13179__A2 _07594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14376__A1 _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16429_ _00817_ clknet_leaf_142_clk register_file\[17\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12926__A2 _07432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10937__A1 _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07802__A1 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11002__I _06220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14679__A2 register_file\[10\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11937__I _06815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09555__A1 _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13351__A2 _07697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10841__I _06115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11362__A1 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10165__A2 register_file\[11\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ _03766_ _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_115_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07995_ _03327_ _03163_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09307__A1 _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ _05030_ _05044_ _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11114__A1 _06290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09665_ _03934_ _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12862__A1 _07395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08530__A2 _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08616_ _03940_ _03941_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09596_ _04876_ _04908_ _04641_ net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14983__I _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08547_ _03790_ _03793_ net4 _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12614__A1 _07230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12090__A2 _06902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08478_ _03801_ _03804_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13599__I _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14367__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12917__A2 _07425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10440_ _05738_ _05739_ _05740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10928__A1 _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10371_ _03897_ _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12110_ _06652_ _06912_ _06920_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13090_ _07539_ register_file\[16\]\[13\] _07540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09546__A1 _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13342__A2 _07697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12041_ _01874_ _06874_ _06879_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10156__A2 register_file\[18\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11353__A1 _06375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15095__A2 register_file\[8\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15800_ _00188_ clknet_leaf_261_clk register_file\[19\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11105__A1 _06290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13992_ _01508_ register_file\[8\]\[4\] _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09849__A2 register_file\[18\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16297__D _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12943_ _07293_ _07439_ _07445_ _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15731_ _00119_ clknet_leaf_177_clk register_file\[27\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12853__A1 _07388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11656__A2 _06630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10700__B _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15662_ _00050_ clknet_leaf_147_clk register_file\[2\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12874_ _07304_ _07398_ _07403_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14613_ _01954_ _02122_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11825_ _06686_ _06744_ _06749_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14893__I _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12605__A1 _07183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15593_ _03090_ register_file\[21\]\[23\] _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14544_ _02032_ _02053_ _02054_ _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11756_ _06703_ _06704_ _06705_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__A1 _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10707_ _05999_ _06002_ _03795_ _06003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14475_ _01038_ _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15967__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11687_ _06650_ register_file\[8\]\[5\] _06657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13426_ _07536_ _07745_ _07748_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16214_ _00602_ clknet_leaf_207_clk register_file\[24\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10638_ _05752_ register_file\[7\]\[30\] _05935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13030__A1 _07300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16145_ _00533_ clknet_leaf_156_clk register_file\[31\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13357_ _07701_ register_file\[29\]\[17\] _07707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09936__B _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10569_ _05865_ _05866_ _05867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10395__A2 register_file\[23\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11592__A1 _06594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12308_ _06978_ _07050_ _07052_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16076_ _00464_ clknet_leaf_251_clk register_file\[4\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13288_ _07558_ _07663_ _07665_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_170_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11757__I _06143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09537__A1 _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15027_ _02527_ _02531_ _02447_ _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12239_ _06995_ register_file\[31\]\[17\] _07005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11895__A2 _06785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_283_clk_I clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13097__A1 _07539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07780_ _03114_ _02945_ _03115_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14833__A2 register_file\[21\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 addrD[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11647__A2 _06623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15929_ _00317_ clknet_leaf_256_clk register_file\[10\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12844__A1 _07274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08287__B _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09450_ _04558_ register_file\[12\]\[12\] _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_298_clk_I clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08401_ _03726_ _03728_ _01170_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09381_ _04558_ register_file\[16\]\[11\] _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08332_ _03652_ _03660_ _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12072__A2 _06895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_221_clk_I clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10083__A1 _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14349__A1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08263_ register_file\[4\]\[29\] _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13021__A1 _07290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08194_ _03522_ _03524_ _03376_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10386__A2 register_file\[15\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11583__A1 _06024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16122__CLK clknet_leaf_253_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11667__I _06639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14043__I _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13324__A2 _07680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11335__A1 _06368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08041__I _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08200__A1 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11886__A2 _06785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08976__I _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07978_ _03310_ _02978_ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09717_ _04219_ _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11638__A2 _06623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09700__A1 _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09648_ _04892_ register_file\[21\]\[15\] _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09579_ _03897_ _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_93_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11610_ _06606_ register_file\[10\]\[9\] _06608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12590_ _07219_ register_file\[22\]\[24\] _07221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11541_ _06402_ _06561_ _06566_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11810__A2 _06737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15001__A2 register_file\[23\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14260_ _01033_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11472_ _06524_ register_file\[12\]\[18\] _06525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13211_ _07582_ _07619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10423_ _05721_ _05722_ _05723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14760__A1 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14191_ register_file\[5\]\[6\] _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12961__I _07455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10377__A2 register_file\[31\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11574__A1 _06436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13142_ _06154_ _07576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10354_ _05587_ register_file\[25\]\[26\] _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09519__A1 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14512__A1 _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13073_ _07527_ register_file\[16\]\[8\] _07528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10285_ _03860_ _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10129__A2 register_file\[8\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11326__A1 _06427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09047__I _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12024_ _06866_ net33 _06869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11877__A2 register_file\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15068__A2 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14815__A2 register_file\[30\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12826__A1 _07374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11629__A2 register_file\[10\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13975_ _01313_ register_file\[19\]\[4\] _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12201__I _06055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15714_ _00102_ clknet_leaf_54_clk register_file\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12926_ _07276_ _07432_ _07435_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14579__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15645_ _00033_ clknet_leaf_302_clk register_file\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12857_ _07388_ register_file\[1\]\[22\] _07394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11808_ _06670_ _06737_ _06739_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08258__A1 _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15576_ _03072_ _02738_ _03073_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12788_ _07298_ _07350_ _07352_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13251__A1 _07638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12054__A2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14527_ register_file\[4\]\[10\] _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11739_ _06691_ _06692_ _06693_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11801__A2 _06730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16145__CLK clknet_leaf_156_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13003__A1 _07477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14458_ _01962_ _01969_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14751__A1 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13409_ _07734_ register_file\[9\]\[5\] _07739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14389_ _01035_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09666__B _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11565__A1 _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10368__A2 register_file\[7\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16128_ _00516_ clknet_leaf_18_clk register_file\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16295__CLK clknet_leaf_80_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_291_clk clknet_5_5__leaf_clk clknet_leaf_291_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_142_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14503__A1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08950_ _04268_ _04271_ _03817_ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13306__A2 _07670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08981__A2 register_file\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16059_ _00447_ clknet_leaf_288_clk register_file\[5\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11317__A1 _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07901_ _01085_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13857__A3 _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08881_ _04061_ register_file\[20\]\[4\] _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11868__A2 _06768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15059__A2 register_file\[27\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12820__B _07372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09930__A1 _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07832_ _03084_ register_file\[26\]\[24\] _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08733__A2 _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14806__A2 register_file\[27\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12817__A1 _07366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09502_ _04750_ register_file\[7\]\[13\] _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12111__I _06913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12293__A2 _07040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09433_ _03867_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_77_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_160_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09364_ _04473_ register_file\[12\]\[11\] _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12045__A2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10056__A1 _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08315_ _01030_ register_file\[8\]\[30\] _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09997__A1 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_40_clk_I clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09295_ _04409_ register_file\[15\]\[10\] _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13793__A2 _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08246_ _03575_ _01188_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08036__I _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_175_clk_I clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15534__A3 _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13877__I _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08177_ _03504_ _03507_ _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_192_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07875__I _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_282_clk clknet_5_4__leaf_clk clknet_leaf_282_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10070_ _05373_ _05374_ _05375_ _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09921__A1 _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16018__CLK clknet_leaf_229_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12808__A1 _07362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13760_ register_file\[3\]\[1\] _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10972_ _06144_ _06206_ _06208_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10295__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12711_ _07232_ register_file\[21\]\[29\] _07305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13691_ _01207_ _01210_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15222__A2 register_file\[17\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12642_ _07254_ _07248_ _07256_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15430_ _02929_ register_file\[9\]\[21\] _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16168__CLK clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12036__A2 _06874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10047__A1 _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15361_ _01147_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09988__A1 _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12573_ _07205_ register_file\[22\]\[17\] _07211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13784__A2 _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11795__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14312_ _01394_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11524_ _06386_ _06554_ _06556_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15292_ _02792_ _02793_ _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14243_ _01325_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09486__B _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11455_ _06510_ register_file\[12\]\[11\] _06515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12691__I _07231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13536__A2 register_file\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11547__A1 _06565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_31__f_clk clknet_3_7_0_clk clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10406_ _05637_ register_file\[2\]\[26\] _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14174_ _01688_ register_file\[12\]\[6\] _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08412__A1 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11386_ _06407_ _06472_ _06473_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13125_ _07562_ _07556_ _07564_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08963__A2 register_file\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10337_ _05508_ register_file\[3\]\[25\] _05639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13056_ _07513_ _07505_ _07515_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10268_ _05567_ _05570_ _04078_ _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09912__A1 _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12007_ _06815_ register_file\[5\]\[28\] _06858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10199_ _04148_ _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13958_ _01035_ _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10286__A1 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09140__A2 register_file\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12909_ _07422_ register_file\[18\]\[10\] _07426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13889_ _01403_ _01406_ _01076_ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15213__A2 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15628_ _00016_ clknet_leaf_135_clk register_file\[30\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12027__A2 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13224__A1 _07574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09240__I _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10038__A1 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15559_ _03015_ _03057_ _02888_ net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10589__A2 register_file\[4\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08100_ _03352_ register_file\[10\]\[27\] _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09080_ _03991_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08651__A1 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15516__A3 _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08031_ _03359_ _03363_ _03279_ _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14724__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput40 new_value[7] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11538__A1 _06400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15685__CLK clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08403__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_264_clk clknet_5_18__leaf_clk clknet_leaf_264_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09982_ _05090_ register_file\[12\]\[20\] _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12106__I _06913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11010__I _06220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08933_ _03967_ register_file\[20\]\[5\] _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09903__A1 _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08864_ _04185_ _04186_ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11710__A1 _06663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10513__A2 register_file\[8\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07815_ _01083_ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08795_ _04114_ _04117_ _04118_ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15452__A2 _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13463__A1 _07727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10277__A1 _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14007__A3 _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09416_ _04728_ _04730_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13215__A1 _07565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10029__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09347_ _04319_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_178_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ _04593_ _04594_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08642__A1 _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14715__A1 _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08229_ _01120_ register_file\[27\]\[29\] _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11529__A1 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11240_ _06371_ register_file\[19\]\[1\] _06374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_255_clk clknet_5_16__leaf_clk clknet_leaf_255_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08945__A2 register_file\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11171_ _06326_ register_file\[13\]\[6\] _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12016__I _06862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output75_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10752__A2 _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10122_ _05424_ _05426_ _05427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13556__B _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14930_ _02103_ register_file\[10\]\[15\] _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10053_ _03778_ _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11701__A1 _06665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10504__A2 register_file\[24\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09370__A2 register_file\[9\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14861_ register_file\[7\]\[14\] _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15443__A2 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16600_ _00988_ clknet_leaf_257_clk register_file\[9\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13812_ _01317_ _01330_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12257__A2 _07012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14792_ _01155_ _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13454__A1 _07763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16531_ _00919_ clknet_leaf_174_clk register_file\[14\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10955_ _06113_ _06192_ _06198_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13743_ _01152_ register_file\[6\]\[1\] _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_21_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16462_ _00850_ clknet_leaf_129_clk register_file\[16\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13206__A1 _07555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12009__A2 register_file\[5\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10886_ _06026_ register_file\[30\]\[28\] _06153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13674_ _01194_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08881__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15413_ _02911_ _02912_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12625_ _06045_ _07244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16393_ _00781_ clknet_leaf_97_clk register_file\[18\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11768__A1 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12556_ _07193_ _07201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15344_ _02764_ register_file\[8\]\[20\] _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08633__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11507_ _06545_ _06546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_145_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12487_ _06997_ _07153_ _07159_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15275_ _02442_ register_file\[14\]\[19\] _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14226_ _01572_ register_file\[16\]\[7\] _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08404__I register_file\[25\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11438_ _06380_ _06496_ _06504_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14850__B _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_246_clk clknet_5_17__leaf_clk clknet_leaf_246_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14157_ _01666_ _01669_ _01671_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08936__A2 register_file\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09944__B _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11369_ _06390_ _06458_ _06463_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11940__A1 _06818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13108_ _07550_ _07544_ _07552_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14088_ _01603_ register_file\[14\]\[5\] _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13039_ _06019_ _07502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12496__A2 register_file\[23\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13693__A1 _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16333__CLK clknet_leaf_142_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08580_ _03784_ _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_78_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13445__A1 _07756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10259__A1 _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09113__A2 register_file\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13996__A2 _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16483__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15198__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08872__A1 _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09201_ _04518_ register_file\[27\]\[9\] _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14945__A1 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11759__A1 _06706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09132_ _04449_ _04450_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09063_ _04378_ _04381_ _04382_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10982__A2 _06170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08014_ _03344_ _03346_ _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15370__A1 _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12184__A1 _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_237_clk clknet_5_20__leaf_clk clknet_leaf_237_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11931__A1 _06767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09965_ _05270_ _05271_ _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08916_ _04237_ register_file\[17\]\[5\] _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12487__A2 _07153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09896_ _05002_ register_file\[17\]\[19\] _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13684__A1 _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09352__A2 register_file\[29\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08847_ _03807_ _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12239__A2 register_file\[31\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08778_ _04017_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13436__A1 _07546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11998__A1 _06851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10740_ _06029_ register_file\[30\]\[1\] _06034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08863__A1 _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15850__CLK clknet_leaf_111_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10670__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13739__A2 register_file\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ _03864_ register_file\[20\]\[31\] _05967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15610__I _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12410_ _06999_ _07112_ _07113_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13390_ _07580_ _07682_ _07725_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08615__A1 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12411__A2 register_file\[24\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12341_ _07068_ register_file\[25\]\[20\] _07072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10422__A1 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10754__I _06044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08091__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13130__I _07519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10973__A2 register_file\[2\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15060_ _02397_ register_file\[26\]\[17\] _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14164__A2 _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12272_ _06147_ _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14011_ _01527_ _01355_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08918__A2 register_file\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_228_clk clknet_5_21__leaf_clk clknet_leaf_228_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11223_ _06319_ register_file\[13\]\[28\] _06362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09040__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11922__A1 _06703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16356__CLK clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15113__A1 _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09591__A2 register_file\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11154_ _06318_ _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_68_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_27__f_clk_I clknet_3_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11585__I _06591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10105_ _05406_ _05409_ _04900_ _05410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11085_ _06278_ _06279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_122_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15962_ _00350_ clknet_leaf_253_clk register_file\[8\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12478__A2 _07153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13675__A1 _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10036_ _05339_ _05341_ _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09343__A2 register_file\[20\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14913_ _02417_ _02418_ _02336_ _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10489__A1 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15893_ _00281_ clknet_leaf_216_clk register_file\[11\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14844_ _02096_ register_file\[9\]\[14\] _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14775_ _02027_ register_file\[15\]\[13\] _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11987_ _06689_ _06840_ _06846_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11989__A1 _06844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16514_ _00902_ clknet_leaf_20_clk register_file\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13726_ _01245_ _01117_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10938_ _06082_ _06185_ _06188_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08854__A1 _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16445_ _00833_ clknet_leaf_304_clk register_file\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13657_ _00999_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_32_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10869_ _06138_ _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08843__B _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12608_ _06317_ _03836_ _07231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12402__A2 _07105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16376_ _00764_ clknet_leaf_240_clk register_file\[1\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13588_ _01108_ register_file\[8\]\[0\] _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15327_ _02576_ register_file\[17\]\[20\] _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12539_ _07190_ register_file\[22\]\[3\] _07191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10964__A2 register_file\[2\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15258_ _02756_ _02759_ _02508_ _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12166__A1 _06708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_219_clk clknet_5_22__leaf_clk clknet_leaf_219_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14209_ _01635_ register_file\[24\]\[7\] _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13902__A2 register_file\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15189_ _02689_ _02690_ _02691_ _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__I _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11913__A1 _06796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15104__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09582__A2 register_file\[20\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15723__CLK clknet_leaf_136_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09750_ _05052_ _05059_ _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09334__A2 register_file\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08701_ _03837_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_171_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09681_ _04984_ _04991_ _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11141__A2 _06307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ _03831_ _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13418__A1 _07742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07896__A2 register_file\[26\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15873__CLK clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08563_ _03889_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13969__A2 register_file\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14630__A3 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08845__A1 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08494_ _03820_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12641__A2 register_file\[21\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14918__A1 _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10652__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16229__CLK clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09115_ _04434_ _04294_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10955__A2 _06192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09046_ _04335_ _04366_ _04298_ net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16379__CLK clknet_leaf_284_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14146__A2 register_file\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12157__A1 _06698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09022__A1 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11904__A1 _06796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09948_ _05254_ register_file\[16\]\[20\] _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09879_ _04917_ register_file\[25\]\[19\] _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11132__A2 _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11910_ _06691_ _06799_ _06800_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13409__A1 _07734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12890_ _07409_ _07414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10891__A1 _06026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11841_ _06755_ register_file\[7\]\[25\] _06759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10749__I _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14560_ _01904_ register_file\[30\]\[11\] _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11772_ _06163_ _06716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08836__A1 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12632__A2 _07248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10723_ _05989_ _06018_ _03935_ net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13511_ _01031_ register_file\[20\]\[0\] _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14491_ _02000_ _02001_ _01919_ _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09759__B _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16230_ _00618_ clknet_leaf_82_clk register_file\[23\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13442_ _07756_ register_file\[9\]\[19\] _07758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10654_ _05949_ _05950_ _05951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16161_ _00549_ clknet_leaf_65_clk register_file\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13373_ _07562_ _07711_ _07716_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10585_ _05881_ _05882_ _05883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10946__A2 _06192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15112_ _02612_ _02615_ _02447_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12324_ _07061_ register_file\[25\]\[13\] _07062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14137__A2 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07811__A2 register_file\[18\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16092_ _00480_ clknet_leaf_301_clk register_file\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12255_ _06125_ _07016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15043_ _01277_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15746__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13896__A1 _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11206_ _06117_ _06351_ _06352_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12186_ _06036_ _06967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11371__A2 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11137_ _06144_ _06307_ _06309_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12204__I _06059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15945_ _00333_ clknet_leaf_41_clk register_file\[8\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11068_ _06266_ _04067_ _06267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11123__A2 _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12320__A1 _06990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10019_ _05192_ register_file\[19\]\[21\] _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15876_ _00264_ clknet_leaf_62_clk register_file\[11\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14827_ _02164_ register_file\[19\]\[14\] _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10882__A1 _06148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14758_ _02244_ _02265_ _01930_ _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13820__A1 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12623__A2 register_file\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10634__A1 _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13709_ _01227_ _01228_ _01076_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_177_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14689_ _02196_ _02112_ _02197_ _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16428_ _00816_ clknet_leaf_140_clk register_file\[17\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15573__A1 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14376__A2 _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12387__A1 _07094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10394__I _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16359_ _00747_ clknet_leaf_82_clk register_file\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10937__A2 register_file\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12139__A1 _06933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07917__B _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11362__A2 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09802_ _05078_ _05111_ _04977_ net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07994_ _03325_ _03326_ _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09733_ _05038_ _05043_ _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11114__A2 register_file\[27\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09664_ _04959_ _04975_ _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12862__A2 register_file\[1\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08615_ _03786_ register_file\[31\]\[1\] _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09595_ _04891_ _04907_ _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16051__CLK clknet_leaf_231_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08818__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08546_ _03869_ _03872_ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15619__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12614__A2 _07233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10625__A1 _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12784__I _07321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08477_ _03803_ register_file\[28\]\[0\] _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09491__A1 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08294__A2 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10518__B _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09243__A1 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08046__A2 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10928__A2 register_file\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11050__A1 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15316__A1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10370_ _05665_ _05670_ _04655_ _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09029_ _04347_ _04349_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12040_ _06878_ net41 _06879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09546__A2 _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11353__A2 _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12550__A1 _06980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13991_ _01107_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11105__A2 register_file\[27\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12302__A1 _06972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15730_ _00118_ clknet_leaf_173_clk register_file\[27\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12942_ _07443_ register_file\[18\]\[24\] _07445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12853__A2 register_file\[1\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15661_ _00049_ clknet_leaf_142_clk register_file\[2\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14055__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12873_ _07359_ register_file\[1\]\[29\] _07403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14612_ register_file\[4\]\[11\] _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11824_ _06748_ register_file\[7\]\[18\] _06749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08809__A1 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12605__A2 register_file\[22\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15592_ _01134_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13802__A1 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16544__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10616__A1 _05909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14543_ _01194_ _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12694__I _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11755_ _06699_ register_file\[8\]\[25\] _06705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__A2 register_file\[19\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15555__A1 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10706_ _06000_ _06001_ _06002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14474_ _01818_ register_file\[28\]\[10\] _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11686_ _06655_ _06656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16213_ _00601_ clknet_leaf_183_clk register_file\[24\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13425_ _07742_ register_file\[9\]\[12\] _07748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10637_ _05750_ register_file\[6\]\[30\] _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13030__A2 _07494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16144_ _00532_ clknet_leaf_156_clk register_file\[31\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11041__A1 _06117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13356_ _07546_ _07704_ _07706_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10568_ _05609_ register_file\[15\]\[29\] _05866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13581__A3 _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12307_ _07046_ register_file\[25\]\[6\] _07052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16075_ _00463_ clknet_leaf_251_clk register_file\[4\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13287_ _07660_ register_file\[14\]\[21\] _07665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10499_ _05666_ register_file\[6\]\[28\] _05798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09537__A2 register_file\[25\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15026_ _02528_ _02529_ _02530_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_29_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12238_ _06103_ _07004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14530__A2 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12541__A1 _07190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12169_ _06911_ register_file\[3\]\[29\] _06955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14294__A1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16074__CLK clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08568__B _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 addrD[4] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15928_ _00316_ clknet_leaf_264_clk register_file\[10\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12844__A2 _07384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10855__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15859_ _00247_ clknet_leaf_176_clk register_file\[12\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08400_ _03727_ _01097_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09380_ _04556_ register_file\[17\]\[11\] _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08331_ _03655_ _03659_ _01394_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10607__A1 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09473__A1 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15911__CLK clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10083__A2 register_file\[24\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08262_ _03589_ _03591_ _03369_ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14349__A2 register_file\[12\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09225__A1 _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08193_ _03523_ _03374_ _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13021__A2 _07487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11032__A1 _06240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12780__A1 _07347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10852__I _06124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12532__A1 _07186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11335__A2 register_file\[19\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16417__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09862__B _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input37_I new_value[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12779__I _07310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14285__A1 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07977_ _03309_ _03225_ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15155__I _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11099__A1 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09716_ _05024_ _05026_ _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16567__CLK clknet_leaf_215_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09700__A2 _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09647_ _04951_ _04958_ _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09578_ _04883_ _04890_ _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12599__A1 _07183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08529_ _03855_ _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09464__A1 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11540_ _06565_ register_file\[11\]\[13\] _06566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09102__B _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11471_ _06494_ _06524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12019__I _06865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09216__A1 _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08941__B _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11023__A1 _06240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13210_ _07560_ _07615_ _07618_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10422_ _05589_ register_file\[20\]\[27\] _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09767__A2 _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14190_ _01531_ _01704_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07778__A1 _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11858__I _06766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12771__A1 _07281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11574__A2 _06582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10762__I _06051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13141_ _07574_ _07568_ _07575_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10353_ _05650_ _05653_ _04323_ _05654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13072_ _07506_ _07527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14512__A2 register_file\[13\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10284_ _05581_ _05585_ _04018_ _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12523__A1 _07135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16097__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12023_ _01268_ _06864_ _06868_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14276__A1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13974_ _01489_ _01490_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12826__A2 register_file\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15713_ _00101_ clknet_leaf_53_clk register_file\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12925_ _07429_ register_file\[18\]\[17\] _07435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15934__CLK clknet_leaf_305_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10002__I _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15644_ _00032_ clknet_leaf_282_clk register_file\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12856_ _07286_ _07391_ _07393_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14579__A2 register_file\[23\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11807_ _06734_ register_file\[7\]\[11\] _06739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15575_ _02903_ register_file\[31\]\[23\] _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12787_ _07347_ register_file\[20\]\[26\] _07352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13251__A2 register_file\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13313__I _07679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09012__B _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11262__A1 _06388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14526_ _02034_ _02036_ _01702_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11738_ _06687_ register_file\[8\]\[20\] _06693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14457_ _01968_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13003__A2 register_file\[17\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11669_ _06643_ register_file\[8\]\[0\] _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11014__A1 _06069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13408_ _07737_ _07738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_190_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14751__A2 register_file\[21\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14388_ _01818_ register_file\[28\]\[9\] _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12762__A1 _07271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11565__A2 _06575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16127_ _00515_ clknet_leaf_18_clk register_file\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13339_ _07529_ _07690_ _07696_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09238__I _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16058_ _00446_ clknet_leaf_248_clk register_file\[5\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11317__A2 _06420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12514__A1 _07023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15009_ _02513_ register_file\[9\]\[16\] _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07900_ _03068_ register_file\[28\]\[25\] _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08880_ _04059_ register_file\[21\]\[4\] _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07831_ _02998_ register_file\[27\]\[24\] _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07941__A1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12817__A2 register_file\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09501_ _04748_ register_file\[6\]\[13\] _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10828__A1 _06104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09694__A1 _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09432_ _04745_ _04746_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14319__I _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09363_ _04471_ register_file\[13\]\[11\] _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10847__I _06120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10056__A2 register_file\[27\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08314_ _03625_ _03642_ _01505_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_162_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09294_ _04407_ register_file\[14\]\[10\] _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09997__A2 register_file\[2\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08245_ _03574_ _01186_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11005__A1 _06050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08176_ _03505_ _03506_ _01025_ _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14742__A2 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12753__A1 _07326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11678__I _06642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15807__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12505__A1 _07164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13893__I _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08185__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07891__I _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14258__A1 _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15957__CLK clknet_leaf_221_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10971_ _06203_ register_file\[2\]\[26\] _06208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12710_ _06155_ _07304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10295__A2 register_file\[9\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11492__A1 _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13690_ _01208_ _01209_ _01026_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12641_ _07255_ register_file\[21\]\[8\] _07256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14430__A1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10047__A2 register_file\[15\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11244__A1 _06375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15360_ _02858_ _02529_ _02860_ _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_12_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12572_ _07002_ _07208_ _07210_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09988__A2 _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14981__A2 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12992__A1 _07262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14311_ _01822_ _01480_ _01823_ _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11795__A2 register_file\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11523_ _06550_ register_file\[11\]\[6\] _06556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_282_clk_I clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15291_ _01021_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_183_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14242_ _01755_ register_file\[22\]\[7\] _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14733__A2 _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11454_ _06395_ _06513_ _06514_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12744__A1 _07326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10405_ _05702_ _05705_ _05037_ _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11385_ _06469_ register_file\[26\]\[15\] _06473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14173_ _01129_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13124_ _07563_ register_file\[16\]\[23\] _07564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15289__A3 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_297_clk_I clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10336_ _05637_ register_file\[2\]\[25\] _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14497__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10267_ _05568_ _05569_ _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13055_ _07514_ register_file\[16\]\[3\] _07515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12006_ _06708_ _06854_ _06857_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09912__A2 register_file\[21\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_220_clk_I clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10198_ _05501_ register_file\[22\]\[23\] _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07923__A1 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13957_ _01387_ register_file\[28\]\[4\] _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12908_ _07417_ _07425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_235_clk_I clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16112__CLK clknet_leaf_226_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13888_ _01405_ register_file\[26\]\[3\] _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15627_ _00015_ clknet_leaf_99_clk register_file\[30\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12839_ _07269_ _07377_ _07383_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09428__A1 _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14421__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13224__A2 _07622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13043__I _07503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10038__A2 register_file\[31\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15558_ _03034_ _03056_ _02886_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08100__A1 _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14509_ _02018_ _02019_ _01859_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12882__I _07406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15489_ _02903_ register_file\[23\]\[22\] _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08030_ _03360_ _03361_ _03362_ _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput30 new_value[27] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 new_value[8] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10616__B _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11538__A2 _06561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09600__A1 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08403__A2 register_file\[24\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09981_ _05088_ register_file\[13\]\[20\] _05288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14602__I _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08932_ _03965_ register_file\[21\]\[5\] _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13160__A1 _07586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09903__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08863_ _03967_ register_file\[24\]\[4\] _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11710__A2 register_file\[8\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07814_ _03068_ register_file\[20\]\[24\] _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08794_ _04001_ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09667__A1 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11474__A1 _06524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09415_ _04729_ register_file\[4\]\[12\] _04730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13215__A2 _07615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11226__A1 _06156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10029__A2 register_file\[7\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09346_ _04661_ register_file\[22\]\[11\] _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08047__I _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12974__A1 _07244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09277_ _04320_ register_file\[7\]\[10\] _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08642__A2 register_file\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08491__B _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08228_ _03557_ _01117_ _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11529__A2 _06554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12726__A1 _07314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08159_ _03486_ _03489_ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11170_ _06050_ _06330_ _06331_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14479__A1 _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10121_ _05425_ register_file\[12\]\[22\] _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output68_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10052_ _05356_ _05357_ _05358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08510__I _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07905__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11701__A2 _06656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12032__I _06873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14860_ _02033_ register_file\[6\]\[14\] _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_76_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16135__CLK clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13811_ _01322_ _01329_ _01237_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14791_ register_file\[3\]\[13\] _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14651__A1 _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11871__I _06769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13454__A2 register_file\[9\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16530_ _00918_ clknet_leaf_175_clk register_file\[14\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11465__A1 _06517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13742_ _01252_ _01261_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10954_ _06196_ register_file\[2\]\[19\] _06198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16461_ _00849_ clknet_5_27__leaf_clk register_file\[16\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13673_ _01193_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16285__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13206__A2 _07615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_191_clk clknet_5_25__leaf_clk clknet_leaf_191_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10885_ _06151_ _06152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08881__A2 register_file\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15412_ _01065_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11217__A1 _06355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12624_ _07241_ _07233_ _07243_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16392_ _00780_ clknet_leaf_82_clk register_file\[18\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14954__A2 _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11768__A2 _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12965__A1 _07230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15343_ _02825_ _02843_ _02762_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12555_ _06985_ _07194_ _07200_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08633__A2 register_file\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07796__I _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11506_ _06542_ _06545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15274_ _02774_ _02609_ _02775_ _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14706__A2 _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12486_ _07157_ register_file\[23\]\[14\] _07159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12717__A1 _07232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14225_ _01731_ _01738_ _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12207__I _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11437_ _06502_ register_file\[12\]\[4\] _06504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14182__A3 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13390__A1 _07580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14156_ _01670_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11368_ _06462_ register_file\[26\]\[8\] _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13107_ _07551_ register_file\[16\]\[18\] _07552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10319_ _05617_ _05620_ _05421_ _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14087_ _01138_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11299_ _06415_ register_file\[19\]\[18\] _06416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09516__I _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13038_ _07308_ _07458_ _07501_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09897__A1 _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14890__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09649__A1 _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_174_clk_I clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14989_ _02159_ register_file\[17\]\[16\] _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14642__A1 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13445__A2 register_file\[9\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11456__A1 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10259__A2 _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_54_clk_I clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08321__A1 _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_182_clk clknet_5_22__leaf_clk clknet_leaf_182_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_179_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08872__A2 register_file\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09200_ _03810_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11208__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_189_clk_I clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15652__CLK clknet_leaf_69_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11759__A2 _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12956__A1 _07306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09131_ _04172_ register_file\[19\]\[8\] _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_69_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09821__A1 _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13501__I _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09062_ _03795_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_112_clk_I clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10346__B _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12708__A1 _07232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16008__CLK clknet_leaf_296_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08013_ _03345_ register_file\[9\]\[26\] _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08388__A1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13381__A1 _07715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10195__A1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_127_clk_I clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09964_ _05004_ register_file\[24\]\[20\] _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15122__A2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16158__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11177__B _06335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08915_ _03799_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10081__B _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09895_ _05199_ _05202_ _04529_ _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08846_ _04167_ _04168_ _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15425__A3 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08777_ _04099_ _04100_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14633__A1 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13436__A2 _07752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_173_clk clknet_5_29__leaf_clk clknet_leaf_173_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_output106_I net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10670_ _03861_ register_file\[21\]\[31\] _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12947__A1 _07443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09329_ _04441_ register_file\[26\]\[11\] _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12340_ _07049_ _07071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09110__B _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08505__I _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08091__A3 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12271_ _07026_ _07024_ _07027_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08379__A1 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13372__A1 _07715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14010_ register_file\[7\]\[4\] _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11222_ _06148_ _06358_ _06361_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10186__A1 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09040__A2 register_file\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11866__I _06769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10770__I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11922__A2 _06806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11153_ _06319_ _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_68_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13124__A1 _07563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10104_ _05407_ _05408_ _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11084_ _06270_ _06278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15961_ _00349_ clknet_leaf_257_clk register_file\[8\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09879__A1 _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10035_ _05340_ register_file\[28\]\[21\] _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14912_ _02252_ register_file\[18\]\[15\] _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15892_ _00280_ clknet_leaf_213_clk register_file\[11\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14843_ _02349_ register_file\[8\]\[14\] _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12697__I _06138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11438__A1 _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14774_ _02025_ register_file\[14\]\[13\] _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11986_ _06844_ register_file\[5\]\[19\] _06846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15675__CLK clknet_leaf_284_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08303__A1 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16513_ _00901_ clknet_leaf_22_clk register_file\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11989__A2 register_file\[5\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13725_ _01244_ _01115_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10937_ _06182_ register_file\[2\]\[12\] _06188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_164_clk clknet_5_31__leaf_clk clknet_leaf_164_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08854__A2 register_file\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16444_ _00832_ clknet_leaf_286_clk register_file\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14927__A2 _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13656_ _01176_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10868_ _06137_ _06138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12938__A1 _07288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12607_ _06020_ _07230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_169_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16375_ _00763_ clknet_leaf_202_clk register_file\[1\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13587_ _01107_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10799_ _06081_ _06082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15326_ _02826_ register_file\[16\]\[20\] _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12538_ _07185_ _07190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11610__A1 _06606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15257_ _02757_ _02592_ _02758_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12469_ _07142_ register_file\[23\]\[7\] _07149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13363__A1 _07553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14208_ _01674_ _01722_ _01634_ net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12166__A2 _06950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16300__CLK clknet_leaf_139_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15188_ _01074_ _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09031__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11776__I _06718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11913__A2 register_file\[6\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14139_ _01644_ _01653_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13115__A1 _07555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13991__I _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16450__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08700_ _04023_ _04024_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09690__B _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09680_ _04987_ _04990_ _04026_ _04991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08542__A1 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08631_ _03956_ register_file\[6\]\[1\] _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13418__A2 register_file\[9\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11429__A1 _06366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08562_ _03783_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14091__A2 _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_155_clk clknet_5_30__leaf_clk clknet_leaf_155_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08493_ _03798_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_165_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08845__A2 register_file\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14918__A2 register_file\[22\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12929__A1 _07278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14327__I _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09114_ _04431_ _04432_ _04433_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11601__A1 _06598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08073__A3 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09045_ _04352_ _04365_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13354__A1 _07543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12157__A2 _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10168__A1 _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09022__A2 register_file\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11686__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11904__A2 register_file\[6\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08781__A1 _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09947_ _03863_ _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09878_ _05182_ _05185_ _04094_ _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15698__CLK clknet_leaf_178_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08829_ _03917_ register_file\[2\]\[3\] _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13409__A2 register_file\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11840_ _06729_ _06758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_166_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10891__A2 register_file\[30\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12093__A1 _06863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_146_clk clknet_5_27__leaf_clk clknet_leaf_146_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11771_ _06714_ _06643_ _06715_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13510_ _01030_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10722_ _06004_ _06017_ _06018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14909__A2 _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14490_ _01835_ register_file\[18\]\[10\] _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13441_ _07550_ _07752_ _07757_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10765__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14237__I _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10653_ _03890_ register_file\[15\]\[30\] _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16160_ _00548_ clknet_leaf_12_clk register_file\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13372_ _07715_ register_file\[29\]\[23\] _07716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10584_ _05695_ register_file\[23\]\[29\] _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15111_ _02613_ _02529_ _02614_ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12323_ _07041_ _07061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16091_ _00479_ clknet_leaf_288_clk register_file\[4\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13345__A1 _07694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15042_ _02546_ _02378_ _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12254_ _07014_ _07012_ _07015_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13896__A2 register_file\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11205_ _06348_ register_file\[13\]\[20\] _06352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16473__CLK clknet_leaf_202_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12185_ _06965_ _06961_ _06966_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08772__A1 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11136_ _06304_ register_file\[27\]\[26\] _06309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11659__A1 _06591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15944_ _00332_ clknet_leaf_44_clk register_file\[8\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11067_ _06265_ _06266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12320__A2 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10018_ _05190_ register_file\[18\]\[21\] _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15017__B _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15875_ _00263_ clknet_leaf_50_clk register_file\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10331__A1 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14826_ _02332_ _02249_ _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10882__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14757_ _02255_ _02264_ _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_137_clk clknet_5_26__leaf_clk clknet_leaf_137_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11969_ _06830_ register_file\[5\]\[12\] _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13708_ _01072_ register_file\[26\]\[1\] _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11831__A1 _06748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14688_ _02027_ register_file\[15\]\[12\] _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16427_ _00815_ clknet_leaf_141_clk register_file\[17\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13639_ _01153_ _01157_ _01159_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15573__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12387__A2 register_file\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16358_ _00746_ clknet_leaf_82_clk register_file\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10398__A1 _05689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09252__A2 _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15309_ _02809_ _01066_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12890__I _07409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16289_ _00677_ clknet_leaf_68_clk register_file\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13336__A1 _07694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10624__B _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11898__A1 _06679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ _05097_ _05110_ _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08763__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15840__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07993_ _02993_ register_file\[25\]\[26\] _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14836__A1 _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09732_ _05042_ _04973_ _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14610__I _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08515__A1 _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09663_ _04966_ _04974_ _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08614_ _03780_ register_file\[30\]\[1\] _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09594_ _04901_ _04906_ _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08545_ _03871_ register_file\[15\]\[0\] _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08818__A2 register_file\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11822__A1 _06684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10625__A2 register_file\[17\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08476_ _03802_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09491__A2 register_file\[23\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15564__A2 _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09243__A2 register_file\[30\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10389__A1 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15316__A2 register_file\[28\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16496__CLK clknet_leaf_174_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11050__A2 _06250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_300_clk clknet_5_4__leaf_clk clknet_leaf_300_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09028_ _04348_ register_file\[27\]\[6\] _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11889__A1 _06782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12550__A2 _07194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14827__A1 _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10561__A1 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13990_ _01484_ _01504_ _01506_ _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output50_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08506__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12302__A2 _07040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12941_ _07290_ _07439_ _07444_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10313__A1 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13136__I _06146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15660_ _00048_ clknet_leaf_135_clk register_file\[2\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12872_ _07302_ _07398_ _07402_ _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15252__A1 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14055__A2 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14611_ _02117_ _02119_ _02120_ _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11823_ _06718_ _06748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12066__A1 _06892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12975__I _07457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15591_ _01132_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08809__A2 register_file\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13802__A2 register_file\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14542_ _02044_ _02052_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11813__A1 _06674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11754_ _06655_ _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _03785_ register_file\[27\]\[31\] _06001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14473_ _01978_ _01983_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11685_ _06642_ _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15713__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16212_ _00600_ clknet_leaf_157_clk register_file\[24\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13424_ _07534_ _07745_ _07747_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13566__A1 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10636_ _05931_ _05932_ _05933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08037__A3 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16143_ _00531_ clknet_leaf_153_clk register_file\[31\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11041__A2 _06250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13355_ _07701_ register_file\[29\]\[16\] _07706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10567_ _05607_ register_file\[14\]\[29\] _05865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13318__A1 _07682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12306_ _06974_ _07050_ _07051_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08993__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16074_ _00462_ clknet_5_5__leaf_clk register_file\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13286_ _07555_ _07663_ _07664_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10498_ _05795_ _05796_ _05797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10444__B _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_14__f_clk clknet_3_3_0_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15025_ _02444_ register_file\[15\]\[16\] _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12237_ _07002_ _07000_ _07003_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12215__I _06975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08745__A1 _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12168_ _06710_ _06950_ _06954_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_11__f_clk_I clknet_3_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10552__A1 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11119_ _06297_ register_file\[27\]\[19\] _06299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12099_ _06913_ _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14294__A2 register_file\[24\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 addrS[0] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15927_ _00315_ clknet_leaf_220_clk register_file\[10\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09170__A1 _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10855__A2 _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16369__CLK clknet_leaf_160_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15858_ _00246_ clknet_leaf_171_clk register_file\[12\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14809_ _02312_ _02315_ _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12057__A1 _06885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15789_ _00177_ clknet_leaf_123_clk register_file\[19\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ _03656_ _03361_ _03658_ _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_162_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09473__A2 register_file\[24\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08261_ _03590_ _01167_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08192_ register_file\[5\]\[28\] _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09225__A2 register_file\[10\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11032__A2 register_file\[28\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13309__A1 _07631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08984__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12780__A2 register_file\[20\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10791__A1 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12532__A2 register_file\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10543__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11964__I _06825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15436__I _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14340__I _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07976_ _03307_ _03308_ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15482__A1 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09715_ _05025_ register_file\[15\]\[16\] _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11099__A2 _06286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12296__A1 _07042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09161__A1 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09646_ _04954_ _04957_ _04139_ _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09577_ _04886_ _04889_ _04017_ _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15736__CLK clknet_leaf_199_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08528_ _03854_ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12599__A2 register_file\[22\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13796__A1 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09464__A2 register_file\[13\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08267__A3 _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08459_ _03785_ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11204__I _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11470_ _06412_ _06520_ _06523_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15886__CLK clknet_leaf_187_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09216__A2 register_file\[22\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10421_ _05587_ register_file\[21\]\[27\] _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12220__A1 _06990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07778__A2 register_file\[14\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12771__A2 _07336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output98_I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13140_ _07504_ register_file\[16\]\[28\] _07575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10352_ _05651_ _05652_ _05653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13071_ _06062_ _07526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10283_ _05582_ _05584_ _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12523__A2 register_file\[23\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12022_ _06866_ net22 _06868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10534__A1 _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15473__A1 _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16511__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13973_ _01009_ _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12287__A1 _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12924_ _07274_ _07432_ _07434_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15712_ _00100_ clknet_leaf_15_clk register_file\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12855_ _07388_ register_file\[1\]\[21\] _07393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15643_ _00031_ clknet_leaf_271_clk register_file\[30\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13787__A1 _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11806_ _06667_ _06737_ _06738_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15574_ _02736_ register_file\[30\]\[23\] _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12786_ _07295_ _07350_ _07351_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14525_ _02035_ _01786_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11262__A2 _06384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11737_ _06655_ _06692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13539__A1 _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14456_ _01966_ _01967_ _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11668_ _06642_ _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13407_ _07729_ _07737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11014__A2 _06229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10619_ _05731_ register_file\[28\]\[30\] _05916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14387_ _01895_ _01898_ _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11599_ _06593_ _06601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_155_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16126_ _00514_ clknet_leaf_33_clk register_file\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12762__A2 _07336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13338_ _07694_ register_file\[29\]\[9\] _07696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08423__I register_file\[23\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10174__B _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10773__A1 _06042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08430__A3 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16041__CLK clknet_leaf_291_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16057_ _00445_ clknet_leaf_242_clk register_file\[5\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13269_ _07538_ _07649_ _07654_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08718__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15008_ _01110_ _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12514__A2 _07174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13711__A1 _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07830_ _03164_ _02912_ _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14267__A2 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16191__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07941__A2 register_file\[14\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15759__CLK clknet_leaf_146_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09143__A1 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09500_ _04811_ _04813_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10828__A2 _06096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09431_ _04473_ register_file\[8\]\[12\] _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09203__B _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09362_ _04657_ _04677_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08313_ _03634_ _03641_ _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09293_ _04608_ _04609_ _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08244_ _03572_ _03573_ _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11959__I _06817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12202__A1 _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11005__A2 _06229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08175_ _03352_ register_file\[10\]\[28\] _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12753__A2 register_file\[20\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10764__A1 _06050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08421__A3 _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08709__A1 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12505__A2 register_file\[23\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13702__A1 _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16534__CLK clknet_leaf_226_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10516__A1 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14258__A2 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07932__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07959_ _03292_ _03210_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10970_ _06139_ _06206_ _06207_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09629_ _04938_ _04940_ _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11492__A2 _06534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12640_ _07234_ _07255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13769__A1 _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12571_ _07205_ register_file\[22\]\[16\] _07210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12441__A1 _07087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11244__A2 _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_50_clk clknet_5_9__leaf_clk clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14310_ _01650_ register_file\[31\]\[8\] _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11522_ _06382_ _06554_ _06555_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12992__A2 _07473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15290_ _02785_ _02791_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14241_ _01089_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16064__CLK clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11453_ _06510_ register_file\[12\]\[10\] _06514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08948__A1 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09339__I _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12744__A2 register_file\[20\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13941__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ _05703_ _05704_ _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14172_ _01680_ _01686_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11384_ _06457_ _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_125_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08412__A3 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13123_ _07503_ _07563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10335_ _03779_ _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14497__A2 register_file\[23\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13054_ _07506_ _07514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10266_ _05503_ register_file\[31\]\[24\] _05569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10507__A1 _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12005_ _06851_ register_file\[5\]\[27\] _06857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10197_ _04145_ _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15446__A1 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14249__A2 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07923__A2 register_file\[23\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11109__I _06278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13956_ _01469_ _01472_ _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12907_ _07257_ _07418_ _07424_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13887_ _01404_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12838_ _07381_ register_file\[1\]\[14\] _07383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15626_ _00014_ clknet_leaf_99_clk register_file\[30\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09428__A2 _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14421__A2 register_file\[8\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12769_ _07278_ _07336_ _07341_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15557_ _03046_ _03055_ _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_41_clk clknet_5_13__leaf_clk clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08100__A2 register_file\[10\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14508_ _01684_ register_file\[10\]\[10\] _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15488_ _02736_ register_file\[22\]\[22\] _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10994__A1 _06033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11779__I _06721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14155__I _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput20 new_value[18] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14439_ register_file\[7\]\[9\] _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput31 new_value[28] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput42 new_value[9] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10746__A1 _06037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16109_ _00497_ clknet_leaf_192_clk register_file\[3\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09980_ _05283_ _05286_ _04057_ _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14488__A2 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08931_ _04249_ _04252_ _03877_ _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12499__A1 _07009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09364__A1 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13160__A2 register_file\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12403__I _07089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08862_ _03965_ register_file\[25\]\[4\] _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15437__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11171__A1 _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07813_ _03144_ _03147_ _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07914__A2 _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08793_ _04115_ _04116_ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09667__A2 register_file\[25\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09712__I _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12671__A1 _07267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10858__I _06129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13234__I _07630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09414_ _03823_ _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08328__I _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14412__A2 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09345_ _04316_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16087__CLK clknet_leaf_234_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12423__A1 _07116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11226__A2 _06358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_32_clk clknet_5_6__leaf_clk clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_179_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12974__A2 _07456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09276_ _04317_ register_file\[6\]\[10\] _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11689__I _06055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08227_ _03556_ _01115_ _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08158_ _03487_ _03488_ _03168_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08089_ _03420_ register_file\[31\]\[27\] _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08998__I _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15924__CLK clknet_leaf_209_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14479__A2 register_file\[31\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10120_ _04415_ _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_99_clk clknet_5_15__leaf_clk clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10051_ _05090_ register_file\[24\]\[21\] _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13151__A2 _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15428__A1 _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07905__A2 register_file\[31\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13853__B _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09107__A1 _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13810_ _01324_ _01326_ _01328_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14790_ _02131_ register_file\[2\]\[13\] _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_5_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14651__A2 register_file\[17\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13741_ _01256_ _01260_ _01148_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12662__A1 _07269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10953_ _06108_ _06192_ _06197_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08330__A2 _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16460_ _00848_ clknet_leaf_131_clk register_file\[16\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13672_ net10 _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10884_ _06150_ _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14403__A2 _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15411_ _02910_ _02746_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12623_ _07242_ register_file\[21\]\[3\] _07243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12414__A1 _07004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16391_ _00779_ clknet_leaf_82_clk register_file\[18\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12983__I _07457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11217__A2 register_file\[13\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_23_clk clknet_5_3__leaf_clk clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15342_ _02835_ _02842_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12554_ _07198_ register_file\[22\]\[9\] _07200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08094__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12965__A2 _07456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10976__A1 _06152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11599__I _06593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11505_ _06543_ _06544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_157_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15273_ _02610_ register_file\[13\]\[19\] _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12485_ _06994_ _07153_ _07158_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14224_ _01734_ _01737_ _01395_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_172_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11436_ _06377_ _06496_ _06503_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09594__A1 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14155_ _01051_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13390__A2 _07682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11367_ _06449_ _06462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13106_ _07503_ _07551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10318_ _05618_ _05619_ _05620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14086_ _01600_ _01343_ _01601_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08701__I _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11298_ _06367_ _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09346__A1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13037_ _07455_ register_file\[17\]\[31\] _07501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10249_ _05418_ register_file\[7\]\[24\] _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15419__A1 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14890__A2 register_file\[27\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13763__B _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09649__A2 register_file\[20\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14988_ _02411_ register_file\[16\]\[16\] _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11456__A2 _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13939_ _01454_ _01456_ _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13054__I _07506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13989__I _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12405__A1 _06994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11208__A2 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15609_ _02936_ register_file\[10\]\[23\] _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16589_ _00977_ clknet_leaf_117_clk register_file\[9\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07987__I _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_14_clk clknet_5_2__leaf_clk clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_50_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09130_ _04170_ register_file\[18\]\[8\] _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08085__A1 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12956__A2 _07410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09821__A2 register_file\[13\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10967__A1 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09061_ _04379_ _04380_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07832__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15947__CLK clknet_leaf_115_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08012_ _01013_ _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09585__A1 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08388__A2 register_file\[14\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13381__A2 register_file\[29\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11392__A1 _06476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10195__A2 register_file\[20\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09963_ _05002_ register_file\[25\]\[20\] _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09337__A1 _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08914_ _04231_ _04235_ _04037_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09894_ _05200_ _05201_ _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11144__A1 _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09888__A2 _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14769__B _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ _03803_ register_file\[16\]\[4\] _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12892__A1 _07241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_281_clk_I clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08776_ _03811_ register_file\[19\]\[3\] _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14633__A2 register_file\[25\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input12_I new_value[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12644__A1 _07255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_296_clk_I clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07897__I _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09328_ _04642_ _04643_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12947__A2 register_file\[18\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08076__A1 _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10958__A1 _06117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14149__A1 _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09259_ _03785_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12270_ _07019_ register_file\[31\]\[26\] _07027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11221_ _06355_ register_file\[13\]\[27\] _06361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13372__A2 register_file\[29\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11383__A1 _06405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10186__A2 register_file\[13\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output80_I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_234_clk_I clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11152_ _06318_ _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08521__I _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10103_ _05275_ register_file\[23\]\[22\] _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13124__A2 register_file\[16\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14321__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15960_ _00348_ clknet_leaf_242_clk register_file\[8\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11083_ _06046_ _06269_ _06277_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11135__A1 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09879__A2 register_file\[25\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14872__A2 _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13675__A3 _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14911_ _02164_ register_file\[19\]\[15\] _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10034_ _03900_ _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_249_clk_I clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15891_ _00279_ clknet_leaf_213_clk register_file\[11\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08677__B _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14842_ _01079_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14624__A2 _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12635__A1 _07250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11438__A2 _06496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14773_ _02279_ _02192_ _02280_ _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11985_ _06686_ _06840_ _06845_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16512_ _00900_ clknet_leaf_1_clk register_file\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10936_ _06078_ _06185_ _06187_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13724_ _01241_ _01243_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14388__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16443_ _00831_ clknet_leaf_274_clk register_file\[17\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10867_ net28 _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13655_ _01175_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13602__I _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12938__A2 _07439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12606_ _07036_ _07186_ _07229_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08067__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13586_ _00993_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16374_ _00762_ clknet_leaf_223_clk register_file\[1\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10949__A1 _06189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10798_ _06080_ _06081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15325_ _01107_ _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07814__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12537_ _06967_ _07184_ _07189_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12218__I _06077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11610__A2 register_file\[10\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12468_ _06978_ _07146_ _07148_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15256_ _02593_ register_file\[31\]\[19\] _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09567__A1 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14560__A1 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13363__A2 _07704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14207_ _01698_ _01721_ _01632_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11419_ _06447_ register_file\[26\]\[30\] _06492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15187_ _02520_ register_file\[10\]\[18\] _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12399_ _07102_ register_file\[24\]\[11\] _07107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11374__A1 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14138_ _01647_ _01652_ _01395_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13115__A2 _07556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09971__B _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14069_ _01323_ register_file\[22\]\[5\] _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11126__A1 _06297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_clk clknet_5_0__leaf_clk clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I addrD[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12874__A1 _07304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11792__I _06729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08630_ _03827_ _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08542__A2 register_file\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08561_ _03887_ register_file\[10\]\[0\] _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11429__A2 _06496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12626__A1 _07242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08492_ _03797_ _03818_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14379__A1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14608__I register_file\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13512__I _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12929__A2 _07432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08058__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13051__A1 _07507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08606__I _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09113_ _04291_ register_file\[1\]\[7\] _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07805__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09044_ _04359_ _04364_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16125__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13668__B _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15343__A3 _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09558__A1 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13354__A2 _07704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10168__A2 register_file\[25\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11365__A1 _06454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08230__A1 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16275__CLK clknet_leaf_209_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08781__A2 register_file\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09946_ _05252_ register_file\[17\]\[20\] _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11117__A1 _06297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14854__A2 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12865__A1 _07395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09877_ _05183_ _05184_ _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09730__A1 _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08828_ _04144_ _04151_ _03914_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _04083_ _03929_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12617__A1 _07237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10111__I _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11770_ _06640_ register_file\[8\]\[30\] _06715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08297__A1 _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13290__A1 _07560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12093__A2 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10721_ _06011_ _06016_ _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15031__A2 _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13440_ _07756_ register_file\[9\]\[18\] _07757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10652_ _03887_ register_file\[14\]\[30\] _05949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09797__A1 _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14790__A1 _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13371_ _07678_ _07715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10583_ _05693_ register_file\[22\]\[29\] _05881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12322_ _06992_ _07057_ _07060_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15110_ _02444_ register_file\[15\]\[17\] _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16090_ _00478_ clknet_leaf_248_clk register_file\[4\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_173_clk_I clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15041_ _02538_ _02545_ _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12253_ _07007_ register_file\[31\]\[21\] _07015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14542__A1 _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10781__I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11356__A1 _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09347__I _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11204_ _06329_ _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_53_clk_I clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12184_ _06963_ register_file\[31\]\[1\] _06966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15098__A2 _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ _06139_ _06307_ _06308_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08772__A2 register_file\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11108__A1 _06091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_188_clk_I clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15642__CLK clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15943_ _00331_ clknet_leaf_43_clk register_file\[8\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11066_ _03783_ net43 _06265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12856__A1 _07286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_68_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10017_ _05321_ _05322_ _05323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09721__A1 _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15874_ _00262_ clknet_leaf_50_clk register_file\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10331__A2 register_file\[30\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_111_clk_I clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14825_ _02330_ _02331_ _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12608__A1 _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15792__CLK clknet_leaf_169_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14756_ _02260_ _02263_ _02091_ _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13281__A1 _07550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12084__A2 _06902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11968_ _06670_ _06833_ _06835_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10095__A1 _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10956__I _06177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13707_ _01069_ register_file\[27\]\[1\] _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10919_ _06169_ _06177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_126_clk_I clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14687_ _02025_ register_file\[14\]\[12\] _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11831__A2 register_file\[7\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11899_ _06789_ register_file\[6\]\[16\] _06794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15022__A2 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16426_ _00814_ clknet_leaf_98_clk register_file\[17\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16148__CLK clknet_leaf_151_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13638_ _01158_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13033__A1 _07455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09788__A1 _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16357_ _00745_ clknet_leaf_74_clk register_file\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13569_ _01089_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10398__A2 _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11595__A1 _06598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15308_ _02807_ _02808_ _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08460__A1 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16288_ _00676_ clknet_leaf_16_clk register_file\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16298__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13336__A2 register_file\[29\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15239_ _02735_ _02740_ _02658_ _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08212__A1 _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11898__A2 _06792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09800_ _05104_ _05109_ _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08763__A2 register_file\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07992_ _03243_ register_file\[24\]\[26\] _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14836__A2 register_file\[23\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13639__A3 _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09731_ _05039_ _05040_ _05041_ _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10640__B _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14112__B _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09662_ _04972_ _04973_ _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08613_ _03937_ _03938_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09593_ _04905_ _04637_ _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11027__I _06228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08544_ _03870_ _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08279__A1 _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10086__A1 _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13811__A3 _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08475_ _03771_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11822__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13242__I _07633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09779__A1 _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14772__A1 _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15169__I _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09027_ _03889_ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11338__A1 _06368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09167__I _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15665__CLK clknet_leaf_173_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13878__A3 _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09951__A1 _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12838__A1 _07381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09929_ _04967_ register_file\[2\]\[19\] _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09703__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08506__A2 register_file\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12940_ _07443_ register_file\[18\]\[23\] _07444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11510__A1 _06546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12871_ _07359_ register_file\[1\]\[28\] _07402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14610_ _01158_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11822_ _06684_ _06744_ _06747_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13263__A1 _07646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15590_ _03003_ register_file\[20\]\[23\] _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12066__A2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10776__I _06062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14541_ _02051_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11753_ _06138_ _06703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11813__A2 _06737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13152__I _07582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10704_ _03916_ register_file\[26\]\[31\] _06000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13015__A1 _07484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14472_ _01979_ _01981_ _01982_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11684_ _06049_ _06654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08690__A1 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16211_ _00599_ clknet_leaf_157_clk register_file\[24\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13423_ _07742_ register_file\[9\]\[11\] _07747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13566__A2 register_file\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10635_ _03844_ register_file\[4\]\[30\] _05932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09786__B _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16440__CLK clknet_leaf_204_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11577__A1 _06543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16142_ _00530_ clknet_leaf_153_clk register_file\[31\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13354_ _07543_ _07704_ _07705_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08442__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10566_ _05862_ _05863_ _05864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12305_ _07046_ register_file\[25\]\[5\] _07051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14515__A1 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08993__A2 register_file\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13318__A2 register_file\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13285_ _07660_ register_file\[14\]\[20\] _07664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16073_ _00461_ clknet_leaf_289_clk register_file\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10497_ _05731_ register_file\[4\]\[28\] _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11329__A1 _06427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12236_ _06995_ register_file\[31\]\[16\] _07003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15024_ _01693_ _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16590__CLK clknet_leaf_188_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09942__A1 _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08745__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12167_ _06911_ register_file\[3\]\[28\] _06954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14818__A2 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09805__I _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10552__A2 register_file\[18\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11118_ _06108_ _06293_ _06298_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12829__A1 _07374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12098_ _06910_ _06913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_110_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13327__I _07681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12231__I _06094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11049_ _06254_ register_file\[28\]\[24\] _06256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15926_ _00314_ clknet_leaf_203_clk register_file\[10\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 addrS[1] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11501__A1 _06495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09170__A2 register_file\[13\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15857_ _00245_ clknet_leaf_171_clk register_file\[12\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14808_ _02313_ _02314_ _01982_ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13254__A1 _07524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12057__A2 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15788_ _00176_ clknet_leaf_123_clk register_file\[19\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09540__I _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10068__A1 _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14739_ _02245_ _02246_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13062__I _07519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08260_ register_file\[7\]\[29\] _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13006__A1 _07276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14754__A1 _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16409_ _00797_ clknet_leaf_263_clk register_file\[18\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08191_ _03203_ _03521_ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10240__A1 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13309__A2 register_file\[14\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08984__A2 register_file\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10791__A2 _06074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13946__B _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14621__I _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10543__A2 register_file\[28\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07975_ _03222_ register_file\[17\]\[26\] _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10370__B _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15482__A2 register_file\[18\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09714_ _03889_ _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09161__A2 register_file\[25\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13681__B _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09645_ _04955_ _04956_ _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09576_ _04887_ _04888_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12048__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13245__A1 _07638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08527_ _03790_ _03793_ net4 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14993__A1 _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13796__A2 register_file\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16463__CLK clknet_leaf_148_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_20__f_clk clknet_3_5_0_clk clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08458_ _03784_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08672__A1 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14745__A1 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08389_ _01015_ register_file\[15\]\[31\] _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11559__A1 _06572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10420_ _05716_ _05719_ _04323_ _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12220__A2 _06988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_285_clk clknet_5_5__leaf_clk clknet_leaf_285_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10351_ _05583_ register_file\[19\]\[26\] _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12316__I _07049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13070_ _07524_ _07520_ _07525_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10282_ _05583_ register_file\[19\]\[25\] _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12021_ _01163_ _06864_ _06867_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13720__A2 _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07854__B _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11731__A1 _06687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09625__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_3__f_clk_I clknet_3_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12051__I _06865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12287__A2 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13972_ _01487_ _01488_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10298__A1 _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15711_ _00099_ clknet_leaf_15_clk register_file\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12923_ _07429_ register_file\[18\]\[16\] _07434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15225__A2 _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08685__B _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15642_ _00030_ clknet_5_18__leaf_clk register_file\[30\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12854_ _07283_ _07391_ _07392_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13236__A1 _07634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11805_ _06734_ register_file\[7\]\[10\] _06738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14984__A1 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15573_ _03069_ _02733_ _03070_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12785_ _07347_ register_file\[20\]\[25\] _07351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11798__A1 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14524_ register_file\[7\]\[10\] _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11736_ _06116_ _06691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08663__A1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10470__A1 _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14455_ _01800_ register_file\[1\]\[9\] _01801_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11667_ _06639_ _06642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13406_ _07516_ _07728_ _07736_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10618_ _05729_ register_file\[29\]\[30\] _05915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08704__I _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14386_ _01896_ _01897_ _01560_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11598_ _06380_ _06592_ _06600_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10455__B _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16125_ _00513_ clknet_leaf_34_clk register_file\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_276_clk clknet_5_7__leaf_clk clknet_leaf_276_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13337_ _07526_ _07690_ _07695_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10549_ _05587_ register_file\[17\]\[29\] _05847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10773__A2 register_file\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11970__A1 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16056_ _00444_ clknet_leaf_244_clk register_file\[5\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13268_ _07653_ register_file\[14\]\[13\] _07654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15537__I register_file\[7\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09915__A1 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15007_ _02349_ register_file\[8\]\[16\] _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08718__A2 register_file\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12219_ _06983_ register_file\[31\]\[11\] _06991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13199_ _07582_ _07612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11722__A1 _06679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16336__CLK clknet_leaf_162_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09391__A2 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08194__A3 _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13057__I _06044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13475__A1 _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09143__A2 register_file\[21\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15909_ _00297_ clknet_leaf_63_clk register_file\[10\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12896__I _07417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16486__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14019__A3 _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09430_ _04471_ register_file\[9\]\[12\] _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13227__A1 _07583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ _04666_ _04676_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14975__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11305__I _06383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11789__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08312_ _03637_ _03640_ _03340_ _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_178_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09292_ _04473_ register_file\[12\]\[10\] _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08654__A1 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10461__A1 _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08243_ _03345_ register_file\[9\]\[29\] _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08174_ _03350_ register_file\[11\]\[28\] _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12202__A2 register_file\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10213__A1 _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_267_clk clknet_5_18__leaf_clk clknet_leaf_267_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_192_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12136__I _06921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13950__A2 _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10764__A2 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11961__A1 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15152__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09906__A1 _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input42_I new_value[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07958_ _03286_ _03291_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13466__A1 _07576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07889_ _03222_ register_file\[25\]\[25\] _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15182__I _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09628_ _04939_ register_file\[11\]\[15\] _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13218__A1 _07567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08893__A1 _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09180__I _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15853__CLK clknet_leaf_126_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14966__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13769__A2 register_file\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09559_ _04870_ _04871_ _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12570_ _06999_ _07208_ _07209_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08645__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12441__A2 register_file\[24\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11521_ _06550_ register_file\[11\]\[5\] _06555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14240_ _01752_ _01410_ _01753_ _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11452_ _06505_ _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15391__A1 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08524__I _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10403_ _05503_ register_file\[11\]\[26\] _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14171_ _01683_ _01685_ _01431_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08948__A2 register_file\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11383_ _06405_ _06465_ _06471_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09070__A1 _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16359__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10334_ _05632_ _05635_ _04139_ _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13122_ _06128_ _07562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13053_ _06039_ _07513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14261__I _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10265_ _05501_ register_file\[30\]\[24\] _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11704__A1 _06663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12004_ _06706_ _06854_ _06856_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10196_ _05498_ _05499_ _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15446__A2 register_file\[15\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14249__A3 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13457__A1 _07763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13955_ _01470_ _01471_ _01026_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13605__I _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12906_ _07422_ register_file\[18\]\[9\] _07424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09304__B _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13209__A1 _07612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08884__A1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13886_ _01029_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15625_ _00013_ clknet_leaf_100_clk register_file\[30\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14957__A1 _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12837_ _07266_ _07377_ _07382_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15556_ _03054_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12768_ _07340_ register_file\[20\]\[18\] _07341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14507_ _01682_ register_file\[11\]\[10\] _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11719_ _06094_ _06679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15487_ _02984_ _02733_ _02985_ _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_187_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13340__I _07689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12699_ _07291_ register_file\[21\]\[25\] _07297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10994__A2 _06219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14438_ _01611_ register_file\[6\]\[9\] _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xinput10 addrS[4] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 new_value[19] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 new_value[29] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10185__B _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput43 we net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_249_clk clknet_5_16__leaf_clk clknet_leaf_249_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_50_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14369_ register_file\[3\]\[8\] _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10746__A2 _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11943__A1 _06645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16108_ _00496_ clknet_leaf_193_clk register_file\[3\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15726__CLK clknet_leaf_146_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08930_ _04250_ _04251_ _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16039_ _00427_ clknet_leaf_296_clk register_file\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12499__A2 _07160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09265__I _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09364__A2 register_file\[12\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08861_ _04179_ _04182_ _04183_ _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11171__A2 register_file\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07812_ _03145_ _03146_ _02814_ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10204__I _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13448__A1 _07558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08792_ _03851_ register_file\[11\]\[3\] _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15876__CLK clknet_leaf_62_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12120__A1 _06926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13515__I _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08609__I _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08875__A1 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12671__A2 register_file\[21\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10682__A1 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09413_ _04727_ register_file\[5\]\[12\] _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09344_ _04658_ _04659_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08627__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12423__A2 register_file\[24\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10434__A1 _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09275_ _04590_ _04591_ _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14346__I _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08226_ _03554_ _03555_ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14176__A2 _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07850__A2 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12187__A1 _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08157_ _01090_ register_file\[18\]\[28\] _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09052__A1 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11934__A1 _06716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08088_ _01096_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09175__I _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10050_ _05088_ register_file\[25\]\[21\] _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15428__A2 register_file\[8\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09107__A2 register_file\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13740_ _01257_ _01258_ _01259_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10952_ _06196_ register_file\[2\]\[18\] _06197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08866__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12662__A2 _07260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14939__A1 _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__A1 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16031__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13671_ _01174_ _01191_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10883_ net31 _06150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15410_ _02908_ _02909_ _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12622_ _07234_ _07242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16390_ _00778_ clknet_leaf_82_clk register_file\[18\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12414__A2 _07112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10425__A1 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15341_ _02838_ _02841_ _02508_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_40_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12553_ _06982_ _07194_ _07199_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09291__A1 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08094__A2 register_file\[8\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10976__A2 _06206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11504_ _06542_ _06543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15272_ _02524_ register_file\[12\]\[19\] _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16181__CLK clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12484_ _07157_ register_file\[23\]\[13\] _07158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07841__A2 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15749__CLK clknet_leaf_69_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14223_ _01735_ _01480_ _01736_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09794__B _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09043__A1 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11435_ _06502_ register_file\[12\]\[3\] _06503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11925__A1 _06803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14154_ _01667_ _01326_ _01668_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11366_ _06388_ _06458_ _06461_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08397__A3 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13105_ _06106_ _07550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10317_ _05418_ register_file\[7\]\[25\] _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11297_ _06107_ _06414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14085_ _01344_ register_file\[13\]\[5\] _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13678__A1 _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09346__A2 register_file\[22\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08149__A3 _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15899__CLK clknet_leaf_265_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10248_ _05416_ register_file\[6\]\[24\] _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13036_ _07306_ _07458_ _07500_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12350__A1 _07075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15419__A2 register_file\[29\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10179_ _04124_ _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14987_ _02483_ _02491_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13335__I _07681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12102__A1 _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13938_ _01455_ _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08857__A1 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10664__A1 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13869_ _01030_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15608_ _02934_ register_file\[11\]\[23\] _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12405__A2 _07105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16588_ _00976_ clknet_5_24__leaf_clk register_file\[9\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16524__CLK clknet_leaf_123_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15539_ _03036_ _03037_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08085__A2 register_file\[29\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10967__A2 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09060_ _04172_ register_file\[27\]\[7\] _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14158__A2 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07832__A2 register_file\[26\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12169__A1 _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08011_ _03181_ register_file\[8\]\[26\] _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11916__A1 _06803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09585__A2 register_file\[23\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15107__A1 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09962_ _05264_ _05267_ _05268_ _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09337__A2 register_file\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08913_ _04232_ _04234_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14330__A2 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09893_ _04998_ register_file\[7\]\[19\] _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12341__A1 _07068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14881__A3 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08844_ _03800_ register_file\[17\]\[4\] _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12892__A2 _07408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10869__I _06138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16054__CLK clknet_leaf_234_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08775_ _03808_ register_file\[18\]\[3\] _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08848__A1 _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12644__A2 register_file\[21\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08312__A3 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15460__I _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10407__A1 _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09327_ _04369_ register_file\[24\]\[11\] _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09273__A1 _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08076__A2 register_file\[25\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10958__A2 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14149__A2 register_file\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11080__A1 _06275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09258_ _04441_ register_file\[30\]\[10\] _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08209_ _03537_ _03538_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09189_ _04369_ register_file\[12\]\[9\] _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11907__A1 _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11220_ _06144_ _06358_ _06360_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11383__A2 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11151_ _06317_ _04219_ _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_136_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output73_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ _05273_ register_file\[22\]\[22\] _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11082_ _06275_ register_file\[27\]\[4\] _06277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12332__A1 _07002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11135__A2 _06307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ _05338_ register_file\[29\]\[21\] _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14910_ _02415_ _02249_ _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15890_ _00278_ clknet_leaf_171_clk register_file\[11\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14841_ _02327_ _02346_ _02347_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14085__A1 _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13155__I _07585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14772_ _02193_ register_file\[13\]\[13\] _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__A1 _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12635__A2 _07248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11984_ _06844_ register_file\[5\]\[18\] _06845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13832__A1 _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16547__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16511_ _00899_ clknet_leaf_2_clk register_file\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13723_ _01242_ register_file\[9\]\[1\] _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10935_ _06182_ register_file\[2\]\[11\] _06187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16442_ _00830_ clknet_5_18__leaf_clk register_file\[17\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14388__A2 register_file\[28\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15585__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13654_ _01024_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10866_ _06135_ _06118_ _06136_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12399__A1 _07102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12605_ _07183_ register_file\[22\]\[31\] _07229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09264__A1 _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16373_ _00761_ clknet_leaf_222_clk register_file\[1\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13585_ _01054_ _01103_ _01105_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_157_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11403__I _06446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10797_ net14 _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10949__A2 register_file\[2\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15324_ _02816_ _02824_ _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12536_ _07186_ register_file\[22\]\[2\] _07189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07814__A2 register_file\[20\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15255_ _02590_ register_file\[30\]\[19\] _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09016__A1 _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12467_ _07142_ register_file\[23\]\[6\] _07148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14206_ _01712_ _01720_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09808__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09567__A2 register_file\[10\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08712__I _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11418_ _06440_ _06486_ _06491_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14560__A2 register_file\[30\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15186_ _02518_ register_file\[11\]\[18\] _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12398_ _06987_ _07105_ _07106_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12571__A1 _07205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11374__A2 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14137_ _01648_ _01480_ _01651_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11349_ _06366_ _06448_ _06451_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14068_ _01582_ _01410_ _01583_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_3_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11126__A2 register_file\[27\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13019_ _07454_ _07491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14863__A3 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12874__A2 _07398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14076__A1 _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13065__I _06054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08560_ _03886_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13823__A1 _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12626__A2 register_file\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10637__A1 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08491_ _03805_ _03813_ _03817_ _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09699__B _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15914__CLK clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_1__f_clk clknet_3_0_0_clk clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14379__A2 register_file\[24\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15040__A3 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09255__A1 _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08058__A2 register_file\[16\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13051__A2 register_file\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09112_ _04154_ register_file\[3\]\[7\] _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11062__A1 _06218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07805__A2 register_file\[16\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09043_ _04363_ _04294_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09007__A1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_309_clk_I clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14551__A2 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12562__A1 _06992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15500__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09945_ _03860_ _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12314__A1 _07054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11117__A2 register_file\[27\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11983__I _06814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15455__I register_file\[4\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09876_ _04913_ register_file\[15\]\[19\] _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12865__A2 register_file\[1\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09730__A2 register_file\[1\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10876__A1 _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08827_ _04147_ _04150_ _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14067__A1 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08758_ _04080_ _04081_ _04082_ _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_45_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13814__A1 _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12617__A2 _07233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10628__A1 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08297__A2 register_file\[24\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08689_ _03780_ register_file\[18\]\[2\] _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13290__A2 _07663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10720_ _06015_ _03928_ _06016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15567__A1 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10548__B _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10651_ _05946_ _05947_ _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11053__A1 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09797__A2 register_file\[1\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13370_ _07560_ _07711_ _07714_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10582_ _05878_ _05879_ _05880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14790__A2 register_file\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12321_ _07054_ register_file\[25\]\[12\] _07060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10800__A1 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14534__I _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15040_ _02540_ _02543_ _02544_ _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12252_ _06121_ _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12553__A1 _06982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11356__A2 _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11203_ _06113_ _06344_ _06350_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12183_ _06032_ _06965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08221__A2 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11134_ _06304_ register_file\[27\]\[25\] _06308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11108__A2 _06286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12305__A1 _07046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07980__A1 _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15942_ _00330_ clknet_leaf_49_clk register_file\[8\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11065_ _06164_ _06221_ _06264_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12856__A2 _07391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10016_ _05254_ register_file\[16\]\[21\] _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09721__A2 register_file\[8\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15873_ _00261_ clknet_leaf_23_clk register_file\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14058__A1 _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15937__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14824_ _01114_ _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12608__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13805__A1 _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10619__A1 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14755_ _02261_ _02175_ _02262_ _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15314__B _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14709__I _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11967_ _06830_ register_file\[5\]\[11\] _06835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13281__A2 _07656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11292__A1 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13706_ _01224_ _01225_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10095__A2 register_file\[30\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09312__B _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10918_ _06046_ _06168_ _06176_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15558__A1 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14686_ _02191_ _02192_ _02194_ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11898_ _06679_ _06792_ _06793_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16425_ _00813_ clknet_leaf_99_clk register_file\[17\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13637_ _01023_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10849_ _06109_ register_file\[30\]\[21\] _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11133__I _06278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11044__A1 _06247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16356_ _00744_ clknet_leaf_74_clk register_file\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09788__A2 register_file\[13\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13568_ _01029_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14781__A2 _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07799__A1 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15307_ _01062_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12792__A1 _07302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12519_ _07135_ register_file\[23\]\[28\] _07178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_280_clk_I clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16287_ _00675_ clknet_leaf_17_clk register_file\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13499_ _01019_ register_file\[18\]\[0\] _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15238_ _02737_ _02738_ _02739_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14533__A2 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15169_ _01132_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08212__A2 register_file\[19\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_295_clk_I clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ _03315_ _03323_ _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09730_ _04970_ register_file\[1\]\[16\] _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09661_ _04636_ _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14049__A1 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11308__I _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08612_ _03773_ register_file\[28\]\[1\] _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09592_ _04902_ _04903_ _04904_ _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15261__A3 _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08543_ _03784_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09476__A1 _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_233_clk_I clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10086__A2 register_file\[27\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11283__A1 _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08617__I _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08474_ _03800_ register_file\[29\]\[0\] _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14221__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11035__A1 _06247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14772__A2 register_file\[13\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12783__A1 _07293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_248_clk_I clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16242__CLK clknet_leaf_156_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09026_ _04346_ register_file\[26\]\[6\] _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12535__A1 _06965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11338__A2 register_file\[19\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09400__A1 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16392__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14288__A1 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14303__B _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09928_ _05232_ _05235_ _05037_ _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12838__A2 register_file\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10849__A1 _06109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09859_ _04148_ _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12870_ _07300_ _07398_ _07401_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11821_ _06741_ register_file\[7\]\[17\] _06747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13263__A2 register_file\[14\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14460__A1 _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14540_ _02049_ _02050_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11752_ _06701_ _06692_ _06702_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15004__A3 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10703_ _05997_ _05998_ _05999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14471_ _01559_ _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13015__A2 register_file\[17\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14212__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11683_ _06652_ _06641_ _06653_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16210_ _00598_ clknet_leaf_155_clk register_file\[24\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11026__A1 _06091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13422_ _07531_ _07745_ _07746_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10634_ _03841_ register_file\[5\]\[30\] _05931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14763__A2 _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12774__A1 _07283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16141_ _00529_ clknet_leaf_140_clk register_file\[31\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10792__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13353_ _07701_ register_file\[29\]\[15\] _07705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08442__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10565_ _05674_ register_file\[12\]\[29\] _05863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12304_ _07049_ _07050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_143_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14515__A2 register_file\[14\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16072_ _00460_ clknet_leaf_295_clk register_file\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13284_ _07641_ _07663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_136_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10496_ _05729_ register_file\[5\]\[28\] _05795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12526__A1 _07036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11329__A2 register_file\[19\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15023_ _02442_ register_file\[14\]\[16\] _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12235_ _06099_ _07002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09942__A2 register_file\[31\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12166_ _06708_ _06950_ _06953_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12512__I _07145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11117_ _06297_ register_file\[27\]\[18\] _06298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12829__A2 register_file\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12097_ _06911_ _06912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09093__I _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15491__A3 _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11048_ _06130_ _06250_ _06255_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15925_ _00313_ clknet_leaf_218_clk register_file\[10\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11128__I _06267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 addrS[2] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10032__I _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15856_ _00244_ clknet_leaf_170_clk register_file\[12\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16115__CLK clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14807_ _01980_ register_file\[26\]\[14\] _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15787_ _00175_ clknet_leaf_131_clk register_file\[19\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09458__A1 _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14439__I register_file\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12999_ _07269_ _07473_ _07479_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14451__A1 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13254__A2 _07642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11265__A1 _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10068__A2 register_file\[3\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14738_ _02159_ register_file\[17\]\[13\] _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08437__I _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_20__f_clk_I clknet_3_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16265__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13006__A2 _07480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14669_ _02174_ _02175_ _02177_ _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14203__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11017__A1 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16408_ _00796_ clknet_leaf_195_clk register_file\[18\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08190_ register_file\[4\]\[28\] _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14754__A2 register_file\[23\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12765__A1 _07333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16339_ _00727_ clknet_leaf_210_clk register_file\[20\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08433__A2 _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10240__A2 register_file\[15\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14506__A2 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12517__A1 _07171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08197__A1 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13190__A1 _07605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09933__A2 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13518__I _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07974_ _03306_ register_file\[16\]\[26\] _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09713_ _05023_ register_file\[14\]\[16\] _05024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09697__A1 _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09644_ _04691_ register_file\[31\]\[15\] _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_172_clk_I clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09575_ _04691_ register_file\[19\]\[14\] _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09449__A1 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13245__A2 register_file\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11256__A1 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08526_ _03849_ _03852_ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_52_clk_I clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14993__A2 register_file\[19\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10098__B _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09887__B _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08457_ _03783_ _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_187_clk_I clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11008__A1 _06225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14745__A2 register_file\[18\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15632__CLK clknet_leaf_165_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08388_ _01031_ register_file\[14\]\[31\] _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12756__A1 _07333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_67_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08424__A2 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_110_clk_I clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10350_ _05452_ register_file\[18\]\[26\] _05651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12508__A1 _07171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09009_ _04257_ register_file\[22\]\[6\] _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15782__CLK clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10281_ _03919_ _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13181__A1 _07598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12020_ _06866_ net11 _06867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13720__A3 _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_125_clk_I clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11731__A2 register_file\[8\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16138__CLK clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14968__B _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15473__A3 _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13971_ _01062_ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09688__A1 _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15710_ _00098_ clknet_5_3__leaf_clk register_file\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12922_ _07271_ _07432_ _07433_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11495__A1 _06495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15641_ _00029_ clknet_leaf_199_clk register_file\[30\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12853_ _07388_ register_file\[1\]\[20\] _07392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14433__A1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13236__A2 register_file\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11804_ _06729_ _06737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11247__A1 _06378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15572_ _02818_ register_file\[29\]\[23\] _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12784_ _07321_ _07350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14984__A2 register_file\[31\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08112__A1 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11798__A2 _06730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14523_ _02033_ register_file\[6\]\[10\] _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11735_ _06689_ _06680_ _06690_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09860__A1 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08663__A2 register_file\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14454_ _01623_ _01963_ _01965_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10470__A2 register_file\[27\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11666_ _06640_ _06641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_122_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12747__A1 _07257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14208__B _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13405_ _07734_ register_file\[9\]\[4\] _07736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10617_ _05906_ _05913_ _05914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14385_ _01557_ register_file\[26\]\[9\] _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12507__I _07134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08415__A2 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11597_ _06598_ register_file\[10\]\[4\] _06600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08206__B _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16124_ _00512_ clknet_leaf_37_clk register_file\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13336_ _07694_ register_file\[29\]\[8\] _07695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10548_ _05842_ _05845_ _04183_ _05846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16055_ _00443_ clknet_leaf_235_clk register_file\[5\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11970__A2 _06833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15161__A2 _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14722__I _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13267_ _07633_ _07653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10479_ _05765_ _05778_ _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08179__A1 _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15006_ _02492_ _02510_ _02347_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13172__A1 _07522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12218_ _06077_ _06990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09915__A2 register_file\[22\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08720__I _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13198_ _07548_ _07608_ _07611_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11722__A2 _06680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12242__I _06959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12149_ _06940_ register_file\[3\]\[20\] _06944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13475__A2 register_file\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15553__I _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15908_ _00296_ clknet_leaf_62_clk register_file\[10\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11486__A1 _06531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14169__I _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15839_ _00227_ clknet_leaf_13_clk register_file\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11238__A1 _06366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09360_ _04671_ _04674_ _04675_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14975__A2 register_file\[27\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15655__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08103__A1 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12986__A1 _07470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11789__A2 register_file\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08311_ _03638_ _01141_ _03639_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_166_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15502__B _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09291_ _04471_ register_file\[13\]\[10\] _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08654__A2 register_file\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08242_ _01030_ register_file\[8\]\[29\] _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10461__A2 register_file\[30\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12738__A1 _07246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08173_ _03503_ _01188_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11321__I _06138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10213__A2 register_file\[16\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11410__A1 _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15152__A2 register_file\[22\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13163__A1 _07590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13248__I _07641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12910__A1 _07259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input35_I new_value[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07957_ _03288_ _03290_ _02960_ _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13466__A2 _07766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11477__A1 _06524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07888_ _01058_ _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15207__A3 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09627_ _03907_ _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13218__A2 _07622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08893__A2 register_file\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11229__A1 _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09558_ _04602_ register_file\[15\]\[14\] _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12977__A1 _07462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08509_ _03835_ _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_19_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09842__A1 _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09489_ _04801_ _04802_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11520_ _06553_ _06554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_141_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09410__B _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12729__A1 _07239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11451_ _06393_ _06506_ _06512_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15391__A2 register_file\[17\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11231__I _06020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10402_ _05501_ register_file\[10\]\[26\] _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11401__A1 _06476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14170_ _01684_ register_file\[10\]\[6\] _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11382_ _06469_ register_file\[26\]\[14\] _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13867__B _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09070__A2 register_file\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13121_ _07560_ _07556_ _07561_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10333_ _05633_ _05634_ _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13052_ _07511_ _07505_ _07512_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10264_ _05564_ _05566_ _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12901__A1 _07414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12003_ _06851_ register_file\[5\]\[26\] _06856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10195_ _05230_ register_file\[20\]\[23\] _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13457__A2 register_file\[9\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11468__A1 _06410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13954_ _01019_ register_file\[26\]\[4\] _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08333__A1 _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15678__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12905_ _07254_ _07418_ _07423_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14406__A1 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13209__A2 register_file\[15\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_194_clk clknet_5_18__leaf_clk clknet_leaf_194_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13885_ _01313_ register_file\[27\]\[3\] _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08884__A2 register_file\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12836_ _07381_ register_file\[1\]\[13\] _07382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15624_ _00012_ clknet_leaf_89_clk register_file\[30\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14957__A2 register_file\[2\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12968__A1 _07458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15555_ _03050_ _03053_ _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12767_ _07310_ _07340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14506_ _02016_ _01855_ _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11640__A1 _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11718_ _06677_ _06668_ _06678_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15486_ _02818_ register_file\[21\]\[22\] _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12698_ _07247_ _07296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_124_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14437_ _01941_ _01948_ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput11 new_value[0] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11649_ _06627_ register_file\[10\]\[25\] _06631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput22 new_value[1] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput33 new_value[2] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16303__CLK clknet_leaf_145_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14368_ _01713_ register_file\[2\]\[8\] _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13777__B _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13932__A3 _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16107_ _00495_ clknet_leaf_193_clk register_file\[3\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11943__A2 _06816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13319_ _07509_ _07680_ _07684_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14299_ _01810_ _01811_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16038_ _00426_ clknet_leaf_309_clk register_file\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13068__I _06058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16453__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08860_ _03816_ _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08572__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07811_ _02812_ register_file\[18\]\[24\] _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08791_ _03848_ register_file\[10\]\[3\] _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14645__A1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13448__A2 _07759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08324__A1 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12120__A2 register_file\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10131__A1 _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_185_clk clknet_5_28__leaf_clk clknet_leaf_185_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09412_ _03820_ _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_168_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10682__A2 register_file\[31\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15070__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12959__A1 _06316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09343_ _04387_ register_file\[20\]\[11\] _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09824__A1 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08627__A2 register_file\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13531__I _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09274_ _04387_ register_file\[4\]\[10\] _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10434__A2 register_file\[10\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08225_ _01111_ register_file\[25\]\[29\] _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11051__I _06228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13384__A1 _07574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08156_ _01120_ register_file\[19\]\[28\] _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10198__A1 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09052__A2 register_file\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15458__I _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11934__A2 _06770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10890__I _06155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08087_ _01123_ register_file\[30\]\[27\] _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15125__A2 _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13687__A2 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11698__A1 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08989_ _04308_ _04309_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12610__I _07232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08315__A1 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10951_ _06166_ _06196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_44_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_176_clk clknet_5_29__leaf_clk clknet_leaf_176_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08866__A2 register_file\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15970__CLK clknet_leaf_314_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11870__A1 _06652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13670_ _01190_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__A2 register_file\[22\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10882_ _06148_ _06140_ _06149_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12621_ _06040_ _07241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15600__A3 _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15340_ _02839_ _02592_ _02840_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12552_ _07198_ register_file\[22\]\[8\] _07199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11622__A1 _06613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10425__A2 register_file\[23\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09291__A2 register_file\[13\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11503_ _06266_ _04001_ _06542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15271_ _02769_ _02772_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12483_ _07137_ _07157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13375__A1 _07565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14222_ _01650_ register_file\[31\]\[7\] _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11434_ _06497_ _06502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10189__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09043__A2 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11896__I _06777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14153_ _01327_ register_file\[23\]\[6\] _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14272__I _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16476__CLK clknet_leaf_282_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_100_clk clknet_5_15__leaf_clk clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11365_ _06454_ register_file\[26\]\[7\] _06461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13127__A1 _07563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13104_ _07548_ _07544_ _07549_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10316_ _05416_ register_file\[6\]\[25\] _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14084_ _01253_ register_file\[12\]\[5\] _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11296_ _06412_ _06408_ _06413_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13678__A2 _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10305__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13035_ _07455_ register_file\[17\]\[30\] _07500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10247_ _05548_ _05549_ _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08554__A1 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12350__A2 register_file\[25\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10178_ _05481_ register_file\[5\]\[23\] _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14986_ _02486_ _02490_ _02242_ _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08306__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_167_clk clknet_5_31__leaf_clk clknet_leaf_167_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13937_ _01095_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08857__A2 register_file\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11861__A1 _06638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10664__A2 register_file\[8\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13868_ _01381_ _01385_ _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12819_ _07366_ register_file\[1\]\[6\] _07372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15607_ _03103_ _03104_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09806__A1 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16587_ _00975_ clknet_leaf_115_clk register_file\[9\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13799_ _01017_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11613__A1 _06606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15538_ _01354_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15469_ _02634_ register_file\[1\]\[21\] _02635_ _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15355__A2 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13366__A1 _07555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12169__A2 register_file\[3\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08010_ _03324_ _03342_ _03179_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11916__A2 register_file\[6\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15107__A2 register_file\[13\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13118__A1 _07558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15843__CLK clknet_leaf_56_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09961_ _03894_ _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14866__A1 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08912_ _04233_ register_file\[11\]\[5\] _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09892_ _04996_ register_file\[6\]\[19\] _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08545__A1 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12341__A2 register_file\[25\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08843_ _04162_ _04165_ _03962_ _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15993__CLK clknet_leaf_243_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08774_ _04096_ _04097_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_158_clk clknet_5_31__leaf_clk clknet_leaf_158_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08848__A2 register_file\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11046__I _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11852__A1 _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16349__CLK clknet_leaf_302_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10885__I _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14397__A3 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15594__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09326_ _04367_ register_file\[25\]\[11\] _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11604__A1 _06386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09257_ _04572_ _04573_ _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16499__CLK clknet_leaf_174_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09895__B _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11080__A2 register_file\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07823__A3 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13357__A1 _07701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08208_ _03222_ register_file\[17\]\[29\] _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09188_ _04367_ register_file\[13\]\[9\] _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15188__I _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11907__A2 _06792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14092__I _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08139_ _01069_ register_file\[27\]\[28\] _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08304__B _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08784__A1 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11150_ _06316_ _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_175_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10591__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10101_ _05404_ _05405_ _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11081_ _06041_ _06269_ _06276_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12332__A2 _07064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output66_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10032_ _03964_ _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15137__B _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10343__A1 _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12340__I _07049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14840_ _01104_ _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14085__A2 register_file\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14771_ _02107_ register_file\[12\]\[13\] _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11983_ _06814_ _06844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08839__A2 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16510_ _00898_ clknet_leaf_305_clk register_file\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13722_ _01110_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10934_ _06073_ _06185_ _06186_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11843__A1 _06755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13653_ _01172_ _01173_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16441_ _00829_ clknet_leaf_201_clk register_file\[17\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10865_ _06131_ register_file\[30\]\[24\] _06136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15716__CLK clknet_leaf_70_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15585__A2 register_file\[19\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12399__A2 register_file\[24\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12604_ _07034_ _07186_ _07228_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_169_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16372_ _00760_ clknet_leaf_209_clk register_file\[1\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08265__I register_file\[5\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13584_ _01104_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_158_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10796_ _06078_ _06074_ _06079_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09264__A2 register_file\[21\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15323_ _02820_ _02823_ _02658_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12535_ _06965_ _07184_ _07188_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15337__A2 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13348__A1 _07701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15254_ _02754_ _02672_ _02755_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12466_ _06974_ _07146_ _07147_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15866__CLK clknet_leaf_255_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09016__A2 register_file\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14216__B _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14205_ _01719_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12020__A1 _06866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11417_ _06447_ register_file\[26\]\[29\] _06491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15185_ _02686_ _02687_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12397_ _07102_ register_file\[24\]\[10\] _07106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09096__I _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08214__B _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08775__A1 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12571__A2 register_file\[22\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14136_ _01650_ register_file\[31\]\[6\] _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11348_ _06450_ register_file\[26\]\[0\] _06451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14848__A1 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14067_ _01411_ register_file\[21\]\[5\] _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11279_ _06400_ _06396_ _06401_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13018_ _07288_ _07487_ _07490_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15273__A1 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14076__A2 register_file\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12087__A1 _06863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14969_ _00994_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08490_ _03816_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11834__A1 _06696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15025__A1 _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15576__A2 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09255__A2 register_file\[29\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09111_ _04288_ register_file\[2\]\[7\] _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14905__I _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13339__A1 _07529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09042_ _04360_ _04361_ _04362_ _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09007__A2 register_file\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12011__A1 _06815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12562__A2 _07201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10573__A1 _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16021__CLK clknet_leaf_238_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09944_ _05246_ _05250_ _03943_ _05251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15500__A2 register_file\[27\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__A1 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12314__A2 register_file\[25\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13511__A1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09875_ _05117_ register_file\[14\]\[19\] _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__A1 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08826_ _04149_ register_file\[7\]\[3\] _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12160__I _06921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10876__A2 register_file\[30\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16171__CLK clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15264__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14067__A2 register_file\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08757_ _03923_ register_file\[1\]\[2\] _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13814__A2 register_file\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15739__CLK clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11825__A1 _06686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15016__A1 _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08688_ _04011_ _04012_ _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_187_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09494__A2 _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14087__I _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output104_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15567__A2 register_file\[26\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11504__I _06542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10650_ _03883_ register_file\[12\]\[30\] _05947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15889__CLK clknet_leaf_171_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09309_ _04492_ register_file\[10\]\[10\] _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12250__A1 _07007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11053__A2 _06257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15319__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10581_ _05758_ register_file\[20\]\[29\] _05879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_303_clk clknet_5_1__leaf_clk clknet_leaf_303_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12320_ _06990_ _07057_ _07059_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10800__A2 register_file\[30\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12335__I _07038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12251_ _07011_ _07012_ _07013_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12002__A1 _06703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11202_ _06348_ register_file\[13\]\[19\] _06350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08757__A1 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12553__A2 _07194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12182_ _06958_ _06961_ _06964_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10564__A1 _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11133_ _06278_ _06307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_123_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12305__A2 register_file\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16514__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07980__A2 register_file\[18\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15941_ _00329_ clknet_5_8__leaf_clk register_file\[8\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11064_ _06218_ register_file\[28\]\[31\] _06264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10316__A1 _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09182__A1 _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10015_ _05252_ register_file\[17\]\[21\] _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15872_ _00260_ clknet_leaf_7_clk register_file\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15255__A1 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14058__A2 register_file\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14823_ _02328_ _02329_ _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12069__A1 _06892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14754_ _02176_ register_file\[23\]\[13\] _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11966_ _06667_ _06833_ _06834_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15007__A1 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13705_ _01065_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10917_ _06174_ register_file\[2\]\[4\] _06176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11292__A2 register_file\[19\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14685_ _02193_ register_file\[13\]\[12\] _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11897_ _06789_ register_file\[6\]\[15\] _06793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16424_ _00812_ clknet_leaf_83_clk register_file\[17\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13636_ _01154_ _01156_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10848_ _06121_ _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09237__A2 _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14230__A2 _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16355_ _00743_ clknet_leaf_58_clk register_file\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11044__A2 register_file\[28\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13567_ _01082_ _01084_ _01087_ _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_158_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10779_ _06065_ register_file\[30\]\[8\] _06066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07799__A2 register_file\[1\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15306_ _02804_ _02806_ _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12518_ _07028_ _07174_ _07177_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12792__A2 _07350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16286_ _00674_ clknet_leaf_27_clk register_file\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13498_ _01018_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12245__I _06112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15237_ _02488_ register_file\[23\]\[19\] _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12449_ _07135_ _07136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15168_ _02586_ register_file\[28\]\[18\] _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10555__A1 _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08879__B _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14119_ _01590_ _01633_ _01634_ net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15099_ _02602_ _02272_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07990_ _03318_ _03322_ _03075_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16194__CLK clknet_leaf_70_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14297__A2 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09660_ _04968_ _04969_ _04971_ _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14049__A2 register_file\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08920__A1 _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08611_ _03767_ register_file\[29\]\[1\] _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09591_ _04633_ register_file\[1\]\[14\] _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13804__I _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15291__I _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11807__A1 _06734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08542_ _03868_ register_file\[14\]\[0\] _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09476__A2 register_file\[27\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12480__A1 _06990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11283__A2 _06396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08473_ _03799_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14221__A2 register_file\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08987__A1 _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12783__A2 _07343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13980__A1 _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09025_ _03886_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12155__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08739__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12535__A2 _07184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16537__CLK clknet_leaf_241_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09400__A2 register_file\[18\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10546__A1 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15466__I register_file\[3\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14370__I _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15485__A1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14288__A2 register_file\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09927_ _05233_ _05234_ _05235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12299__A1 _07046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09164__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10849__A2 register_file\[30\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _05166_ register_file\[26\]\[18\] _05167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15237__A1 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08809_ _04059_ register_file\[29\]\[3\] _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09789_ _04894_ register_file\[12\]\[17\] _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11820_ _06682_ _06744_ _06746_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11751_ _06699_ register_file\[8\]\[24\] _06702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11234__I _06368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_80_clk clknet_5_11__leaf_clk clknet_leaf_80_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _05758_ register_file\[24\]\[31\] _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14470_ _01980_ register_file\[26\]\[10\] _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11682_ _06650_ register_file\[8\]\[4\] _06653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14212__A2 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13421_ _07742_ register_file\[9\]\[10\] _07746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12223__A1 _06992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11026__A2 _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16067__CLK clknet_leaf_310_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10633_ _05914_ _05929_ _05930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14545__I _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16140_ _00528_ clknet_leaf_139_clk register_file\[31\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08978__A1 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12774__A2 _07343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13352_ _07689_ _07704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10564_ _05672_ register_file\[13\]\[29\] _05862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10785__A1 _06069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12303_ _07041_ _07049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_10_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16071_ _00459_ clknet_leaf_295_clk register_file\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13283_ _07553_ _07656_ _07662_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10495_ _05786_ _05793_ _05794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15022_ _02525_ _02192_ _02526_ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12234_ _06999_ _07000_ _07001_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12526__A2 _07138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13723__A1 _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15376__I _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12165_ _06947_ register_file\[3\]\[27\] _06953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15476__A1 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11116_ _06267_ _06297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12096_ _06910_ _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__A1 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11047_ _06254_ register_file\[28\]\[23\] _06255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15924_ _00312_ clknet_leaf_209_clk register_file\[10\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 addrS[3] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15855_ _00243_ clknet_leaf_127_clk register_file\[12\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14806_ _02230_ register_file\[27\]\[14\] _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15786_ _00174_ clknet_leaf_103_clk register_file\[19\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09458__A2 register_file\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12998_ _07477_ register_file\[17\]\[14\] _07479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14451__A2 register_file\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14737_ _01994_ register_file\[16\]\[13\] _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12462__A1 _06972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11949_ _06822_ register_file\[5\]\[4\] _06824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_71_clk clknet_5_10__leaf_clk clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14668_ _02176_ register_file\[23\]\[12\] _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15400__A1 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14203__A2 register_file\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16407_ _00795_ clknet_leaf_201_clk register_file\[18\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11017__A2 _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13619_ _01139_ register_file\[14\]\[0\] _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14599_ _01776_ register_file\[13\]\[11\] _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12765__A2 register_file\[20\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13962__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16338_ _00726_ clknet_leaf_162_clk register_file\[20\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08453__I _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16269_ _00657_ clknet_leaf_139_clk register_file\[22\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12517__A2 register_file\[23\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13714__A1 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10528__A1 _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09394__A1 _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07944__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07973_ _01055_ _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09146__A1 _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09712_ _03886_ _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09697__A2 register_file\[31\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09643_ _04689_ register_file\[30\]\[15\] _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13534__I _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ _04689_ register_file\[18\]\[14\] _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09449__A2 register_file\[13\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10379__B _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08525_ _03851_ register_file\[19\]\[0\] _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11256__A2 _06384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12453__A1 _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_62_clk clknet_5_9__leaf_clk clknet_leaf_62_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ _03782_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12205__A1 _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11008__A2 register_file\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10893__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07880__A1 _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08387_ _03713_ _01036_ _03714_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13953__A1 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09008_ _04326_ _04328_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12508__A2 register_file\[23\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10280_ _05452_ register_file\[18\]\[25\] _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10519__A1 _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08188__A2 _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13181__A2 register_file\[15\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09137__A1 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14130__A1 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13970_ _01485_ _01486_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09688__A2 register_file\[7\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09922__I _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12921_ _07429_ register_file\[18\]\[15\] _07433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12692__A1 _07291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13444__I _07737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15640_ _00028_ clknet_leaf_197_clk register_file\[30\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12852_ _07369_ _07391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_92_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14433__A2 register_file\[14\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11803_ _06665_ _06730_ _06736_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12783_ _07293_ _07343_ _07349_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15571_ _03068_ register_file\[28\]\[23\] _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12444__A1 _07034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11247__A2 register_file\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_53_clk clknet_5_8__leaf_clk clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11734_ _06687_ register_file\[8\]\[19\] _06690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14522_ _01151_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09860__A2 register_file\[27\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14453_ _01964_ _01883_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14275__I register_file\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11665_ _06639_ _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12747__A2 _07322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13404_ _07513_ _07728_ _07735_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10616_ _05909_ _05912_ _04131_ _05913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14384_ _01813_ register_file\[27\]\[9\] _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11596_ _06377_ _06592_ _06599_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13335_ _07681_ _07694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16123_ _00511_ clknet_leaf_288_clk register_file\[3\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10547_ _05843_ _05844_ _05845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13266_ _07536_ _07649_ _07652_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16054_ _00442_ clknet_leaf_234_clk register_file\[5\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10478_ _05772_ _05777_ _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09376__A1 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12217_ _06987_ _06988_ _06989_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15005_ _02501_ _02509_ _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13172__A2 _07594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13197_ _07605_ register_file\[15\]\[17\] _07611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11183__A1 _06334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12148_ _06921_ _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10930__A1 _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09128__A1 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14121__A1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12079_ _03204_ _06895_ _06901_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15907_ _00295_ clknet_leaf_50_clk register_file\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12683__A1 _07283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_247_clk_I clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16232__CLK clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15838_ _00226_ clknet_leaf_8_clk register_file\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14424__A2 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14894__B _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12435__A1 _07123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11238__A2 _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15769_ _00157_ clknet_leaf_259_clk register_file\[13\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_44_clk clknet_5_12__leaf_clk clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_178_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08103__A2 register_file\[12\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ _03420_ register_file\[31\]\[30\] _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12986__A2 register_file\[17\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09290_ _04589_ _04606_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16382__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08241_ _03553_ _03570_ _01505_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_162_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14185__I register_file\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12738__A2 _07322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13935__A1 _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08172_ _03502_ _01186_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08406__A3 _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11410__A2 _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08911__I _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09367__A1 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09228__B _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11174__A1 _06060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12910__A2 _07425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09119__A1 _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10921__A1 _06174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14112__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07956_ _03289_ _02958_ _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14663__A2 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input28_I new_value[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10888__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07887_ _02889_ register_file\[24\]\[25\] _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09626_ _04937_ register_file\[10\]\[15\] _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14415__A2 _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12426__A1 _07016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09557_ _04600_ register_file\[14\]\[14\] _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14966__A3 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_35_clk clknet_5_6__leaf_clk clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08508_ _03792_ net5 _03793_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_180_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12977__A2 register_file\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09488_ _04669_ register_file\[20\]\[13\] _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08439_ _03765_ _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14095__I _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07853__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11450_ _06510_ register_file\[12\]\[9\] _06512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12729__A2 _07312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10401_ _05700_ _05701_ _05702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11381_ _06402_ _06465_ _06470_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13120_ _07551_ register_file\[16\]\[22\] _07561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output96_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16105__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10332_ _05503_ register_file\[31\]\[25\] _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08821__I _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13439__I _07726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13051_ _07507_ register_file\[16\]\[2\] _07512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10263_ _05565_ register_file\[28\]\[24\] _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11165__A1 _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12002_ _06703_ _06854_ _06855_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12901__A2 register_file\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10194_ _05228_ register_file\[21\]\[23\] _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10912__A1 _06170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08977__B _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16255__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07881__B _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14654__A2 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12665__A1 _07267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11468__A2 _06520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13953_ _01382_ register_file\[27\]\[4\] _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09530__A1 _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12904_ _07422_ register_file\[18\]\[8\] _07423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13884_ _01401_ _01225_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14406__A2 register_file\[18\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15623_ _00011_ clknet_leaf_88_clk register_file\[30\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12417__A1 _07006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12835_ _07361_ _07381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15554_ _03051_ register_file\[1\]\[22\] _03052_ _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_187_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12766_ _07276_ _07336_ _07339_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13090__A1 _07539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10979__A1 _06167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14505_ _02015_ _01853_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11717_ _06675_ register_file\[8\]\[14\] _06678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15485_ _02651_ register_file\[20\]\[22\] _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11640__A2 _06623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12697_ _06138_ _07295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13917__A1 _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14436_ _01944_ _01947_ _01608_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11648_ _06601_ _06630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 new_value[10] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput23 new_value[20] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09597__A1 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput34 new_value[30] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14367_ _01879_ _01538_ _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11579_ _06543_ register_file\[11\]\[30\] _06588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16106_ _00494_ clknet_leaf_41_clk register_file\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13318_ _07682_ register_file\[29\]\[1\] _07684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14298_ _01187_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_171_clk_I clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16037_ _00425_ clknet_leaf_314_clk register_file\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13249_ _07638_ register_file\[14\]\[5\] _07643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11156__A1 _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10903__A1 _06024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07810_ _03063_ register_file\[19\]\[24\] _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08790_ _04112_ _04113_ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_186_clk_I clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14645__A2 register_file\[31\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_66_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09411_ _04718_ _04725_ _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14948__A3 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15772__CLK clknet_leaf_279_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_17_clk clknet_5_2__leaf_clk clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09342_ _04385_ register_file\[21\]\[11\] _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09511__B _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12959__A2 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13081__A1 _07531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09273_ _04385_ register_file\[5\]\[10\] _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_124_clk_I clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08224_ _03243_ register_file\[24\]\[29\] _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16128__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15373__A3 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13384__A2 _07718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08155_ _03485_ _01010_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11395__A1 _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08641__I _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_139_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08086_ _03416_ _03089_ _03417_ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_162_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16278__CLK clknet_leaf_207_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11147__A1 _06164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_19_clk_I clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11698__A2 _06656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09760__A1 _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08988_ _04172_ register_file\[31\]\[6\] _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14636__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07939_ _03271_ _03026_ _03272_ _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11507__I _06545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09512__A1 _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08315__A2 register_file\[8\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10950_ _06104_ _06192_ _06195_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08088__I _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09609_ _04918_ _04920_ _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10881_ _06131_ register_file\[30\]\[27\] _06149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11870__A2 _06768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13722__I _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12620_ _07239_ _07233_ _07240_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_169_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12551_ _07185_ _07198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07826__A1 _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11622__A2 register_file\[10\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11242__I _06036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11502_ _06444_ _06498_ _06541_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12482_ _06992_ _07153_ _07156_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15270_ _02770_ _02771_ _02691_ _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14572__A1 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13375__A2 _07711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14221_ _01478_ register_file\[30\]\[7\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11433_ _06375_ _06496_ _06501_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11386__A1 _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10189__A2 register_file\[14\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14152_ _01323_ register_file\[22\]\[6\] _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11364_ _06386_ _06458_ _06460_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08251__A1 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13127__A2 register_file\[16\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13103_ _07539_ register_file\[16\]\[17\] _07549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10315_ _05615_ _05616_ _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14083_ _01595_ _01598_ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11295_ _06403_ register_file\[19\]\[17\] _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11138__A1 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14875__A2 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15645__CLK clknet_leaf_302_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13678__A3 _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13034_ _07304_ _07494_ _07499_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10246_ _05483_ register_file\[4\]\[24\] _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12886__A1 _07410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12801__I _07359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10177_ _03840_ _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12638__A1 _07252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14985_ _02487_ _02323_ _02489_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15795__CLK clknet_leaf_172_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13936_ register_file\[3\]\[3\] _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11310__A1 _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15333__B _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11861__A2 _06768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13867_ _01383_ _01384_ _01026_ _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15606_ _01426_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12818_ _07246_ _07370_ _07371_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13063__A1 _07514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16586_ _00974_ clknet_leaf_115_clk register_file\[9\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09806__A2 register_file\[20\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13798_ _01312_ _01316_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12248__I _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15537_ register_file\[7\]\[22\] _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12749_ _07326_ register_file\[20\]\[10\] _07330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11613__A2 register_file\[10\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11152__I _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15468_ _02877_ _02965_ _02967_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13366__A2 _07711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14419_ _01910_ _01929_ _01930_ _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__16420__CLK clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15399_ _02651_ register_file\[20\]\[21\] _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11377__A1 _06462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__A1 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13079__I _07519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13118__A2 _07556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14315__A1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09990__A1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _05265_ _05266_ _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11129__A1 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_6_clk clknet_5_0__leaf_clk clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08911_ _03785_ _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16570__CLK clknet_leaf_253_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09891_ _05197_ _05198_ _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12877__A1 _07359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13807__I _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08545__A2 register_file\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ _04163_ _04164_ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08773_ _03803_ register_file\[16\]\[3\] _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11852__A2 _06722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13542__I _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08636__I _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09325_ _04607_ _04640_ _04641_ net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11604__A2 _06602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09256_ _04369_ register_file\[28\]\[10\] _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08207_ _03306_ register_file\[16\]\[29\] _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14554__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09187_ _04470_ _04505_ _04298_ net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11368__A1 _06462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09467__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15668__CLK clknet_leaf_210_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08138_ _03468_ _01066_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08233__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14306__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09981__A1 _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08069_ _03399_ _03150_ _03400_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10100_ _05340_ register_file\[20\]\[22\] _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14857__A2 _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10591__A2 register_file\[6\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11080_ _06275_ register_file\[27\]\[3\] _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12868__A1 _07298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13717__I _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10031_ _05331_ _05336_ _04655_ _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12621__I _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11540__A1 _06565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14609__A2 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_26__f_clk clknet_3_6_0_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_output59_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15282__A2 _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13293__A1 _07562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14770_ _02273_ _02277_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11982_ _06684_ _06840_ _06843_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13721_ _01108_ register_file\[8\]\[1\] _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10933_ _06182_ register_file\[2\]\[10\] _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11843__A2 register_file\[7\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16440_ _00828_ clknet_leaf_204_clk register_file\[17\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10864_ _06134_ _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13045__A1 _07507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13652_ _01051_ _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12603_ _07183_ register_file\[22\]\[30\] _07228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16371_ _00759_ clknet_leaf_211_clk register_file\[1\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12068__I _06873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10795_ _06065_ register_file\[30\]\[11\] _06079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13583_ net10 _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08990__B _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15322_ _02821_ _02738_ _02822_ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12534_ _07186_ register_file\[22\]\[1\] _07188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15253_ _02673_ register_file\[29\]\[19\] _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14283__I register_file\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12465_ _07142_ register_file\[23\]\[5\] _07147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14204_ _01717_ _01718_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13899__A3 _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11416_ _06438_ _06486_ _06490_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08224__A1 _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12396_ _07097_ _07105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15184_ _01426_ _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16593__CLK clknet_leaf_178_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12020__A2 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10031__A1 _05331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14135_ _01649_ _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11347_ _06449_ _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08775__A2 register_file\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11278_ _06391_ register_file\[19\]\[12\] _06401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14066_ _01319_ register_file\[20\]\[5\] _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09724__A1 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13627__I _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13017_ _07484_ register_file\[17\]\[22\] _07490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12531__I _07185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10229_ _05395_ register_file\[9\]\[24\] _05532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13520__A2 _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11531__A1 _06393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_14__f_clk_I clknet_3_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15273__A2 register_file\[13\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14968_ _02429_ _02472_ _02473_ net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12087__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13919_ _01139_ register_file\[14\]\[3\] _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11834__A2 _06751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14899_ _02402_ _02318_ _02404_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13036__A1 _07306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14784__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16569_ _00957_ clknet_leaf_263_clk register_file\[29\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09110_ _04426_ _04429_ _04078_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11598__A1 _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15810__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09041_ _04291_ register_file\[1\]\[6\] _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10270__A1 _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13339__A2 _07690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09963__A1 _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11770__A1 _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10573__A2 register_file\[25\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09943_ _05247_ _05249_ _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13537__I _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09715__A1 _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__A2 register_file\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09236__B _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09874_ _05180_ _05181_ _05182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11522__A1 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16316__CLK clknet_leaf_278_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__A2 register_file\[14\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08825_ _04148_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13275__A1 _07653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12078__A2 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08756_ _03920_ register_file\[3\]\[2\] _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input10_I addrS[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11825__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16466__CLK clknet_leaf_166_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08687_ _03773_ register_file\[16\]\[2\] _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13272__I _07641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13027__A1 _07491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14775__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13578__A2 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11589__A1 _06366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09308_ _04623_ _04624_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10580_ _05756_ register_file\[21\]\[29\] _05878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08454__A1 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12250__A2 register_file\[31\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10261__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _04556_ register_file\[29\]\[9\] _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11520__I _06553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12250_ _07007_ register_file\[31\]\[20\] _07013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08206__A1 _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12002__A2 _06854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11201_ _06108_ _06344_ _06349_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12181_ _06963_ register_file\[31\]\[0\] _06964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11761__A1 _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11132_ _06135_ _06300_ _06306_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09706__A1 _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15940_ _00328_ clknet_leaf_58_clk register_file\[8\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11063_ _06160_ _06221_ _06263_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11513__A1 _06375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10014_ _05316_ _05319_ _03838_ _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09182__A2 register_file\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15871_ _00259_ clknet_leaf_10_clk register_file\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14822_ _02159_ register_file\[17\]\[14\] _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13266__A1 _07536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14753_ _02173_ register_file\[22\]\[13\] _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11965_ _06830_ register_file\[5\]\[10\] _06834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15007__A2 register_file\[8\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13704_ _01223_ _01063_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13018__A1 _07288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10916_ _06041_ _06168_ _06175_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14684_ _01047_ _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11896_ _06777_ _06792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15558__A3 _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15833__CLK clknet_leaf_263_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16423_ _00811_ clknet_leaf_81_clk register_file\[17\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14766__A1 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13635_ _01155_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15611__B _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10847_ _06120_ _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16354_ _00742_ clknet_leaf_58_clk register_file\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13566_ _01086_ register_file\[29\]\[0\] _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10778_ _06028_ _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15305_ _02805_ register_file\[25\]\[20\] _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10252__A1 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12517_ _07171_ register_file\[23\]\[27\] _07177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16285_ _00673_ clknet_leaf_30_clk register_file\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13497_ _01017_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15983__CLK clknet_leaf_245_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15236_ _01325_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15191__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12448_ _07134_ _07135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10004__A1 _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15167_ _02665_ _02669_ _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14741__I _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12379_ _07094_ register_file\[24\]\[3\] _07095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11752__A1 _06701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16339__CLK clknet_leaf_210_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14118_ _01200_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_158_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15098_ _02601_ _02270_ _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14049_ _01564_ register_file\[29\]\[5\] _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input2_I addrD[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15246__A2 _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08920__A2 register_file\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_230_clk clknet_5_21__leaf_clk clknet_leaf_230_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08610_ _03859_ _03932_ _03936_ net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09590_ _04837_ register_file\[3\]\[14\] _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13257__A1 _07526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08541_ _03867_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11807__A2 register_file\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13009__A1 _07278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08472_ _03798_ _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_91_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12480__A2 _07153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10491__A1 _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08987__A2 register_file\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_297_clk clknet_5_4__leaf_clk clknet_leaf_297_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13980__A2 register_file\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11340__I _06163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09024_ _04343_ _04344_ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11991__A1 _06844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08739__A2 register_file\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10546__A2 register_file\[31\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13267__I _07633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15485__A2 register_file\[20\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09926_ _05168_ register_file\[11\]\[19\] _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12299__A2 register_file\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09857_ _04145_ _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15237__A2 register_file\[23\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_221_clk clknet_5_20__leaf_clk clknet_leaf_221_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08808_ _04127_ _04130_ _04131_ _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09788_ _04892_ register_file\[13\]\[17\] _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _03986_ register_file\[26\]\[2\] _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11750_ _06134_ _06701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14748__A1 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10701_ _05756_ register_file\[25\]\[31\] _05997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10482__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11681_ _06045_ _06652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13420_ _07737_ _07745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08824__I _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10632_ _05921_ _05928_ _05929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12223__A2 _06988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_288_clk clknet_5_5__leaf_clk clknet_leaf_288_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13351_ _07541_ _07697_ _07703_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10563_ _05857_ _05860_ _04201_ _05861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10785__A2 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11982__A1 _06684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12302_ _06972_ _07040_ _07048_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15173__A1 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16070_ _00458_ clknet_leaf_309_clk register_file\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13282_ _07660_ register_file\[14\]\[19\] _07662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10494_ _05789_ _05792_ _04262_ _05793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15021_ _02193_ register_file\[13\]\[16\] _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12233_ _06995_ register_file\[31\]\[15\] _07001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14561__I _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13723__A2 register_file\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09655__I _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11734__A1 _06687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12164_ _06706_ _06950_ _06952_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11115_ _06104_ _06293_ _06296_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15476__A2 register_file\[17\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14279__A3 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12095_ _06266_ _03927_ _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__A2 register_file\[8\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11046_ _06217_ _06254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15923_ _00311_ clknet_leaf_213_clk register_file\[10\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_212_clk clknet_5_23__leaf_clk clknet_leaf_212_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13905__I _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09604__B _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15854_ _00242_ clknet_leaf_126_clk register_file\[12\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13239__A1 _07509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14805_ _02311_ _02228_ _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15785_ _00173_ clknet_leaf_103_clk register_file\[19\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12997_ _07266_ _07473_ _07478_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11425__I _06495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14736_ _02234_ _02243_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11948_ _06649_ _06816_ _06823_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12462__A2 _07136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10473__A1 _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14667_ _01096_ _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11879_ _06769_ _06782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13640__I _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15400__A2 register_file\[21\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16406_ _00794_ clknet_leaf_214_clk register_file\[18\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13618_ _01138_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_158_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08734__I _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13411__A1 _07734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14598_ _02107_ register_file\[12\]\[11\] _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10225__A1 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_279_clk clknet_5_6__leaf_clk clknet_leaf_279_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16337_ _00725_ clknet_leaf_157_clk register_file\[20\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13549_ _01069_ register_file\[27\]\[0\] _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13962__A2 register_file\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11973__A1 _06674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16161__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16268_ _00656_ clknet_leaf_138_clk register_file\[22\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15729__CLK clknet_leaf_166_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15219_ _02701_ _02721_ _02471_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14471__I _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14911__A1 _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16199_ _00587_ clknet_leaf_92_clk register_file\[24\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11725__A1 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15467__A2 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07972_ _03261_ _03304_ _03305_ net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15879__CLK clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09146__A2 register_file\[22\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09711_ _05020_ _05021_ _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12150__A1 _06691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_203_clk clknet_5_22__leaf_clk clknet_leaf_203_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09642_ _04952_ _04953_ _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14690__A3 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09573_ _04884_ _04885_ _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08524_ _03850_ _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08657__A1 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12453__A2 _07136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08455_ net1 net2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08386_ _01015_ register_file\[13\]\[31\] _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12205__A2 register_file\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10216__A1 _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13953__A2 register_file\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11070__I _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09909__A1 _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09007_ _04327_ register_file\[20\]\[6\] _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10519__A2 register_file\[29\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13469__A1 _07727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09909_ _05084_ register_file\[31\]\[19\] _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14130__A2 register_file\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11954__B _06827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12141__A1 _06933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12920_ _07417_ _07432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_86_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12692__A2 register_file\[21\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12851_ _07281_ _07384_ _07390_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16034__CLK clknet_leaf_314_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11245__I _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11802_ _06734_ register_file\[7\]\[9\] _06736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15570_ _01080_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12782_ _07347_ register_file\[20\]\[24\] _07349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12444__A2 _07090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14521_ _02021_ _02031_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10455__A1 _05749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11733_ _06112_ _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14452_ register_file\[3\]\[9\] _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__16184__CLK clknet_leaf_191_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11664_ _06216_ _03893_ _06639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13403_ _07734_ register_file\[9\]\[3\] _07735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10615_ _05910_ _05911_ _05912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14383_ _01894_ _01811_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09073__A1 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13944__A2 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11595_ _06598_ register_file\[10\]\[3\] _06599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11955__A1 _06822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16122_ _00510_ clknet_leaf_253_clk register_file\[3\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13334_ _07524_ _07690_ _07693_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10546_ _05583_ register_file\[31\]\[29\] _05844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15387__I _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16053_ _00441_ clknet_leaf_233_clk register_file\[5\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13265_ _07646_ register_file\[14\]\[12\] _07652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10477_ _05776_ _05643_ _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11707__A1 _06663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15004_ _02504_ _02507_ _02508_ _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12216_ _06983_ register_file\[31\]\[10\] _06989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13196_ _07546_ _07608_ _07610_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11183__A2 register_file\[13\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12380__A1 _06969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12147_ _06689_ _06936_ _06942_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10930__A2 register_file\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09128__A2 register_file\[16\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14121__A2 register_file\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12078_ _06899_ net27 _06901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12132__A1 _06933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13635__I _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14672__A3 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11029_ _06095_ _06243_ _06244_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15906_ _00294_ clknet_5_9__leaf_clk register_file\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08729__I _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12683__A2 _07284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13880__A1 _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10694__A1 _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15837_ _00225_ clknet_leaf_279_clk register_file\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11155__I _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15768_ _00156_ clknet_leaf_259_clk register_file\[13\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12435__A2 register_file\[24\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13632__A1 _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16527__CLK clknet_leaf_126_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10446__A1 _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14719_ _02226_ _01976_ _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15699_ _00087_ clknet_leaf_179_clk register_file\[28\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ _03562_ _03569_ _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08464__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12199__A1 _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08171_ _03500_ _03501_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13935__A2 register_file\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15137__A1 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput100 net100 rS[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_133_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11174__A2 _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_7__f_clk clknet_3_1_0_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10921__A2 register_file\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__A2 register_file\[29\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14112__A2 register_file\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07955_ register_file\[5\]\[25\] _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12123__A1 _06665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13545__I _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08639__I _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07886_ _03180_ _03220_ _02888_ net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13871__A1 _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09625_ _03904_ _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_95_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10685__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09556_ _04867_ _04868_ _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12426__A2 _07119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13623__A1 _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08507_ _03829_ _03833_ _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09487_ _04667_ register_file\[21\]\[13\] _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08438_ _03764_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_24_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13926__A2 _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08369_ _03694_ _03695_ _03696_ _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10400_ _05565_ register_file\[8\]\[26\] _05701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11380_ _06469_ register_file\[26\]\[13\] _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08802__A1 _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10331_ _05501_ register_file\[30\]\[25\] _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_307_clk_I clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output89_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13050_ _06035_ _07511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10262_ _03882_ _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14351__A2 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12362__A1 _07032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11165__A2 register_file\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12001_ _06851_ register_file\[5\]\[25\] _06855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10193_ _05489_ _05496_ _05497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08030__A2 _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15300__A1 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14103__A2 _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12114__A1 _06654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08549__I _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13952_ _01467_ _01468_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12665__A2 register_file\[21\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14995__B _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12903_ _07409_ _07422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13883_ _01400_ _01063_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15622_ _00010_ clknet_leaf_89_clk register_file\[30\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12834_ _07264_ _07377_ _07380_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12417__A2 _07112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14286__I _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15553_ _01187_ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12765_ _07333_ register_file\[20\]\[17\] _07339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09294__A1 _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08097__A2 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11703__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10979__A2 register_file\[2\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14504_ _02013_ _02014_ _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11716_ _06090_ _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15484_ _02979_ _02982_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12696_ _07293_ _07284_ _07294_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14435_ _01945_ _01694_ _01946_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_187_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11647_ _06429_ _06623_ _06629_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13917__A2 register_file\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput13 new_value[11] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11928__A1 _06710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09597__A2 register_file\[25\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput24 new_value[21] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14590__A2 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14366_ _01873_ _01878_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput35 new_value[31] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11578_ _06440_ _06582_ _06587_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14235__B _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16105_ _00493_ clknet_leaf_41_clk register_file\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13317_ _07502_ _07680_ _07683_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10529_ _05826_ _05827_ _05828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14297_ _01809_ _01553_ _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16036_ _00424_ clknet_leaf_314_clk register_file\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13248_ _07641_ _07642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12353__A1 _07075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13179_ _07529_ _07594_ _07600_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10903__A2 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10989__I _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12105__A1 _06647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08459__I _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13853__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10667__A1 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09410_ _04721_ _04724_ _03817_ _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09341_ _04648_ _04656_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13081__A2 _07532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09272_ _04579_ _04588_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08223_ _03545_ _03552_ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11919__A1 _06701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08154_ _03484_ _03163_ _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11395__A2 _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08085_ _03090_ register_file\[29\]\[27\] _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14333__A2 _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12344__A1 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11147__A2 _06271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input40_I new_value[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09753__I _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_293_clk_I clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09760__A2 register_file\[21\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08987_ _04170_ register_file\[30\]\[6\] _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07938_ _03027_ register_file\[13\]\[25\] _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09512__A2 _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10658__A1 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07869_ register_file\[4\]\[24\] _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09608_ _04919_ register_file\[16\]\[15\] _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10880_ _06147_ _06148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09539_ _04850_ _04851_ _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09276__A1 _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08079__A2 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_231_clk_I clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11083__A1 _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12550_ _06980_ _07194_ _07197_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15349__A1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07826__A2 register_file\[25\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11501_ _06495_ register_file\[12\]\[31\] _06541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09028__A1 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12481_ _07150_ register_file\[23\]\[12\] _07156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14220_ _01732_ _01475_ _01733_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11432_ _06498_ register_file\[12\]\[2\] _06501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14572__A2 register_file\[18\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_246_clk_I clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12583__A1 _07212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11386__A2 _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14151_ _01664_ _01410_ _01665_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__16222__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09149__B _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11363_ _06454_ register_file\[26\]\[6\] _06460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13102_ _06102_ _07548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10314_ _05483_ register_file\[4\]\[25\] _05616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14082_ _01596_ _01597_ _01431_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_153_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11294_ _06103_ _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11138__A2 register_file\[27\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13033_ _07455_ register_file\[17\]\[29\] _07499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08003__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10245_ _05481_ register_file\[5\]\[24\] _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16372__CLK clknet_leaf_209_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10176_ _05464_ _05479_ _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10897__A1 _06160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14088__A1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14984_ _02488_ register_file\[31\]\[16\] _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12638__A2 _07248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10649__A1 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13935_ _01278_ register_file\[2\]\[3\] _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_35_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11310__A2 _06420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13913__I _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13866_ _01019_ register_file\[18\]\[3\] _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15052__A3 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15605_ _03101_ _03102_ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12817_ _07366_ register_file\[1\]\[5\] _07371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16585_ _00973_ clknet_leaf_114_clk register_file\[9\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12529__I _07183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13063__A2 register_file\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13797_ _01314_ _01315_ _01076_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15536_ _02865_ register_file\[6\]\[22\] _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11074__A1 _06021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12748_ _07321_ _07329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07817__A2 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14744__I _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15467_ _02966_ _02715_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09019__A1 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12679_ _07281_ _07272_ _07282_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14418_ _01505_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14563__A2 _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08742__I _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15398_ _02894_ _02897_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12574__A1 _07004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14349_ _01688_ register_file\[12\]\[8\] _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__A2 register_file\[8\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14315__A2 register_file\[16\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15512__A1 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09990__A2 register_file\[20\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12326__A1 _07061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11129__A2 register_file\[27\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08898__B _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08910_ _04090_ register_file\[10\]\[5\] _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16019_ _00407_ clknet_leaf_228_clk register_file\[6\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09890_ _05063_ register_file\[4\]\[19\] _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08841_ _03786_ register_file\[7\]\[4\] _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14618__A3 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08772_ _03800_ register_file\[17\]\[3\] _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13826__A1 _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15524__B _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08917__I _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09258__A1 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14251__A1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09324_ _03935_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_40_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11065__A1 _06164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07808__A2 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10812__A1 _06091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09255_ _04367_ register_file\[29\]\[10\] _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08206_ _03499_ _03536_ _03305_ net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_154_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09186_ _04488_ _04504_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12565__A1 _06994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08137_ _03467_ _03225_ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09430__A1 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08233__A2 register_file\[28\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16395__CLK clknet_leaf_139_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14306__A2 register_file\[28\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09981__A2 register_file\[13\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08068_ _03235_ register_file\[21\]\[27\] _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12317__A1 _07054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07992__A1 _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12868__A2 _07398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10030_ _05333_ _05335_ _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13817__A1 _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14829__I _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09497__A1 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11981_ _06837_ register_file\[5\]\[17\] _06843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14490__A1 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13293__A2 _07663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13733__I _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13720_ _01220_ _01239_ _01105_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10932_ _06177_ _06185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_147_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_170_clk_I clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13651_ _01160_ _01171_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09249__A1 _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10863_ _06133_ _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14242__A1 _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11253__I _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13045__A2 register_file\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12602_ _07032_ _07222_ _07227_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11056__A1 _06254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16370_ _00758_ clknet_leaf_159_clk register_file\[1\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14793__A2 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_50_clk_I clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13582_ _01078_ _01102_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13889__B _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10794_ _06077_ _06078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15321_ _02488_ register_file\[31\]\[20\] _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12533_ _06958_ _07184_ _07187_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_185_clk_I clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09658__I _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15252_ _02586_ register_file\[28\]\[19\] _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08562__I _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12464_ _07145_ _07146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14203_ _01369_ register_file\[1\]\[6\] _01371_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_65_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11415_ _06447_ register_file\[26\]\[28\] _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15183_ _02684_ _02685_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12395_ _06985_ _07098_ _07104_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09421__A1 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08224__A2 register_file\[24\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14134_ _01095_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11346_ _06446_ _06449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09972__A2 _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12308__A1 _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13908__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07983__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15762__CLK clknet_leaf_177_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14065_ _01577_ _01580_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11277_ _06081_ _06400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13016_ _07286_ _07487_ _07489_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10228_ _05521_ _05530_ _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08527__A3 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11531__A2 _06554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_123_clk_I clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10159_ _05459_ _05462_ _04452_ _05463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16118__CLK clknet_leaf_238_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09488__A1 _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14967_ _01200_ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11295__A1 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13918_ _01434_ _01343_ _01435_ _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_14898_ _02403_ register_file\[29\]\[15\] _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_138_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16268__CLK clknet_leaf_138_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12259__I _06959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13849_ _01177_ _01365_ _01367_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14233__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13036__A2 _07458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11047__A1 _06254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_18_clk_I clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14784__A2 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16568_ _00956_ clknet_leaf_262_clk register_file\[29\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12795__A1 _07311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11598__A2 _06592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15519_ _03016_ _03017_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16499_ _00887_ clknet_leaf_174_clk register_file\[15\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09040_ _04154_ register_file\[3\]\[6\] _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_5_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12547__A1 _07190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09963__A2 register_file\[25\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07974__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11770__A2 register_file\[8\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09942_ _05248_ register_file\[31\]\[20\] _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12722__I _07310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09873_ _05114_ register_file\[12\]\[19\] _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11522__A2 _06554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08824_ _03783_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08755_ _03917_ register_file\[2\]\[2\] _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11286__A1 _06405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08686_ _03767_ register_file\[17\]\[2\] _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08151__A1 _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11038__A1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15635__CLK clknet_leaf_178_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09307_ _04558_ register_file\[8\]\[10\] _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12786__A1 _07295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11589__A2 _06592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09651__A1 _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08454__A2 register_file\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09238_ _03897_ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10261__A2 register_file\[29\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09169_ _04479_ _04487_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11200_ _06348_ register_file\[13\]\[18\] _06349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11210__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12180_ _06962_ _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07965__A1 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11131_ _06304_ register_file\[27\]\[24\] _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11761__A2 register_file\[8\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09427__B _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output71_I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09706__A2 register_file\[19\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11062_ _06218_ register_file\[28\]\[30\] _06263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11513__A2 _06544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10013_ _05317_ _05318_ _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15870_ _00258_ clknet_5_3__leaf_clk register_file\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09941__I _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_6__f_clk_I clknet_3_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14821_ _01994_ register_file\[16\]\[14\] _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14463__A1 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13266__A2 _07649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14752_ _02256_ _02257_ _02259_ _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_166_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11964_ _06825_ _06833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13703_ _01221_ _01222_ _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10915_ _06174_ register_file\[2\]\[3\] _06175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14683_ _01774_ _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13018__A2 _07487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14215__A1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09890__A1 _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11895_ _06677_ _06785_ _06791_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11029__A1 _06095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16422_ _00810_ clknet_leaf_83_clk register_file\[17\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13634_ _01095_ _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10846_ net24 _06120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12777__A1 _07340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16353_ _00741_ clknet_leaf_58_clk register_file\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13565_ _01085_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10777_ _06063_ _06064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15304_ _01058_ _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12516_ _07026_ _07174_ _07176_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14518__A2 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10252__A2 register_file\[25\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16284_ _00672_ clknet_5_6__leaf_clk register_file\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13496_ _00992_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15235_ _02736_ register_file\[22\]\[19\] _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12447_ _06265_ _03991_ _07134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11201__A1 _06108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10004__A2 _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15166_ _02666_ _02668_ _02336_ _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12378_ _07089_ _07094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13741__A3 _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13638__I _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14117_ _01610_ _01631_ _01632_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11752__A2 _06692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11329_ _06427_ register_file\[19\]\[27\] _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15097_ _02599_ _02600_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14048_ _01038_ _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14469__I _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10997__I _06220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13257__A2 _07642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14454__A1 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16090__CLK clknet_leaf_248_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15999_ _00387_ clknet_leaf_0_clk register_file\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11268__A1 _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08540_ _03806_ _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15658__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08133__A1 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ _03764_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__13009__A2 _07480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14206__A1 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10491__A2 register_file\[22\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12768__A1 _07340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09633__A1 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08436__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10243__A2 _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09023_ _04061_ register_file\[24\]\[6\] _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11991__A2 register_file\[5\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13193__A1 _07605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12940__A1 _07443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13548__I _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09925_ _05166_ register_file\[10\]\[19\] _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16433__CLK clknet_leaf_162_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09856_ _05163_ _05164_ _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08807_ _03795_ _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09787_ _05087_ _05096_ _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11259__A1 _06386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08738_ _04060_ _04062_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16583__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08669_ _03898_ register_file\[9\]\[1\] _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09872__A1 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10700_ _05992_ _05995_ _03914_ _05996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11680_ _06649_ _06641_ _06651_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10482__A2 register_file\[16\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12759__A1 _07269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10631_ _05924_ _05927_ _04553_ _05928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15003__I _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13350_ _07701_ register_file\[29\]\[14\] _07703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11431__A1 _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10562_ _05858_ _05859_ _05860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12301_ _07046_ register_file\[25\]\[4\] _07048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11982__A2 _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13281_ _07550_ _07656_ _07661_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14842__I _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10493_ _05790_ _05791_ _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15020_ _02524_ register_file\[12\]\[16\] _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13184__A1 _07534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12232_ _06975_ _07000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14920__A2 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07938__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12931__A1 _07281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12163_ _06947_ register_file\[3\]\[26\] _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11114_ _06290_ register_file\[27\]\[17\] _06296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12094_ _03686_ _06866_ _06909_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15922_ _00310_ clknet_leaf_185_clk register_file\[10\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11045_ _06126_ _06250_ _06253_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11498__A1 _06440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15800__CLK clknet_leaf_261_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15853_ _00241_ clknet_leaf_126_clk register_file\[12\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13239__A2 _07632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11706__I _06077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14804_ _02310_ _01976_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12996_ _07477_ register_file\[17\]\[13\] _07478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15784_ _00172_ clknet_leaf_108_clk register_file\[19\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12998__A1 _07477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14735_ _02238_ _02241_ _02242_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11947_ _06822_ register_file\[5\]\[3\] _06823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09863__A1 _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15950__CLK clknet_leaf_189_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14666_ _01325_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11670__A1 _06638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10473__A2 register_file\[2\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11878_ _06660_ _06778_ _06781_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13617_ _01029_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16405_ _00793_ clknet_leaf_213_clk register_file\[18\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10829_ net20 _06106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09615__A1 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14597_ _01129_ _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13411__A2 register_file\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10225__A2 register_file\[23\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11422__A1 _06444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16306__CLK clknet_leaf_158_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16336_ _00724_ clknet_leaf_162_clk register_file\[20\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13548_ _01068_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_185_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11973__A2 _06833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16267_ _00655_ clknet_leaf_138_clk register_file\[22\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13479_ _00999_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15218_ _02712_ _02720_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16198_ _00586_ clknet_leaf_91_clk register_file\[24\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07929__A1 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12922__A1 _07271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11725__A2 _06680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15149_ _02651_ register_file\[20\]\[18\] _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12272__I _06147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07971_ _01199_ _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09710_ _04756_ register_file\[12\]\[16\] _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11489__A1 _06531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09581__I _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08354__A1 _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12150__A2 _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09641_ _04756_ register_file\[28\]\[15\] _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15219__A3 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14427__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10161__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09572_ _04756_ register_file\[16\]\[14\] _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12989__A1 _07470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08523_ _03784_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_64_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09854__A1 _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09530__B _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11661__A1 _06591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08454_ _03780_ register_file\[26\]\[0\] _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10676__B _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09606__A1 _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08385_ _01031_ register_file\[12\]\[31\] _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08409__A2 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10216__A2 register_file\[19\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11413__A1 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09082__A2 _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09006_ _03843_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13166__A1 _07516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09909__A2 register_file\[31\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08660__I _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14902__A2 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12913__A1 _07422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15823__CLK clknet_leaf_127_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09908_ _05082_ register_file\[30\]\[19\] _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12141__A2 register_file\[3\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09839_ _04124_ _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_24_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15973__CLK clknet_leaf_313_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12850_ _07388_ register_file\[1\]\[19\] _07390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11801_ _06662_ _06730_ _06735_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12781_ _07290_ _07343_ _07348_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08648__A2 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14520_ _02024_ _02029_ _02030_ _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11732_ _06686_ _06680_ _06688_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16329__CLK clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11652__A1 _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10586__B _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14451_ _01713_ register_file\[2\]\[9\] _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11663_ _06020_ _06638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15394__A2 _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13402_ _07729_ _07734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11404__A1 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10207__A2 _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10614_ _03871_ register_file\[27\]\[30\] _05911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14382_ _01893_ _01553_ _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11594_ _06593_ _06598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16121_ _00509_ clknet_leaf_241_clk register_file\[3\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13333_ _07686_ register_file\[29\]\[7\] _07693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10545_ _03828_ register_file\[30\]\[29\] _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_130_clk clknet_5_26__leaf_clk clknet_leaf_130_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13157__A1 _07502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16052_ _00440_ clknet_leaf_230_clk register_file\[5\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13264_ _07534_ _07649_ _07651_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10476_ _05773_ _05774_ _05775_ _05776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_170_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12904__A1 _07422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15003_ _01670_ _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11707__A2 register_file\[8\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12215_ _06975_ _06988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_155_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13195_ _07605_ register_file\[15\]\[16\] _07610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12380__A2 _07088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12146_ _06940_ register_file\[3\]\[19\] _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14657__A1 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12077_ _03123_ _06895_ _06900_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11028_ _06240_ register_file\[28\]\[15\] _06244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15905_ _00293_ clknet_leaf_23_clk register_file\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_197_clk clknet_5_19__leaf_clk clknet_leaf_197_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08887__A2 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13880__A2 register_file\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15836_ _00224_ clknet_leaf_279_clk register_file\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12979_ _07462_ register_file\[17\]\[6\] _07468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15767_ _00155_ clknet_leaf_224_clk register_file\[13\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14718_ _02224_ _02225_ _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09350__B _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15698_ _00086_ clknet_leaf_178_clk register_file\[28\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14649_ _01994_ register_file\[16\]\[12\] _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14188__A3 _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07862__A3 _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12199__A2 register_file\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13396__A1 _07730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08170_ _03345_ register_file\[9\]\[28\] _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16319_ _00707_ clknet_leaf_15_clk register_file\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_121_clk clknet_5_24__leaf_clk clknet_leaf_121_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput101 net101 rS[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__14896__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14360__A3 _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08575__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10382__A1 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15996__CLK clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12730__I _07313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07954_ _03203_ _03287_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08327__A1 _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12123__A2 _06922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13320__A1 _07682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_188_clk clknet_5_25__leaf_clk clknet_leaf_188_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07885_ _03198_ _03219_ _02886_ _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11346__I _06446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13871__A2 register_file\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09624_ _04934_ _04935_ _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11882__A1 _06782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15073__A1 _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09555_ _04669_ register_file\[12\]\[14\] _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14820__A1 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13623__A2 register_file\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08506_ _03832_ register_file\[23\]\[0\] _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11634__A1 _06620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09486_ _04796_ _04799_ _04102_ _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12177__I _06959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08437_ _03763_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_71_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13387__A1 _07679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08368_ _03459_ register_file\[1\]\[31\] _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_149_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09055__A2 _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14392__I _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15128__A2 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_112_clk clknet_5_13__leaf_clk clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08802__A2 register_file\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08299_ _03626_ _03627_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10330_ _05630_ _05631_ _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10261_ _05563_ register_file\[29\]\[24\] _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12000_ _06825_ _06854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_106_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12362__A2 _07078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10192_ _05492_ _05495_ _03876_ _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16001__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12640__I _07234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12114__A2 _06922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13311__A1 _06316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13951_ _01370_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_179_clk clknet_5_23__leaf_clk clknet_leaf_179_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13862__A2 _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12902_ _07252_ _07418_ _07421_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13882_ _01398_ _01399_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15064__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16151__CLK clknet_leaf_190_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12833_ _07374_ register_file\[1\]\[12\] _07380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15621_ _00009_ clknet_leaf_72_clk register_file\[30\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15719__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13471__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11625__A1 _06613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10428__A2 _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12764_ _07274_ _07336_ _07338_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15552_ _01004_ _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09294__A2 register_file\[14\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14503_ _01676_ register_file\[9\]\[10\] _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11715_ _06674_ _06668_ _06676_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15483_ _02980_ _02981_ _02814_ _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12695_ _07291_ register_file\[21\]\[24\] _07294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15367__A2 _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13378__A1 _07567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14434_ _01605_ register_file\[15\]\[9\] _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11646_ _06627_ register_file\[10\]\[24\] _06629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 new_value[12] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11928__A2 _06806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12815__I _07361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14365_ _01875_ _01877_ _01709_ _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput25 new_value[22] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_103_clk clknet_5_15__leaf_clk clknet_leaf_103_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput36 new_value[3] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11577_ _06543_ register_file\[11\]\[29\] _06587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16104_ _00492_ clknet_leaf_42_clk register_file\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13316_ _07682_ register_file\[29\]\[0\] _07683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07909__I _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10600__A2 _05897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10528_ _05565_ register_file\[12\]\[28\] _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14296_ _01807_ _01808_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13247_ _07633_ _07641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16035_ _00423_ clknet_leaf_314_clk register_file\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10335__I _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10459_ _05758_ register_file\[28\]\[27\] _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08557__A1 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13178_ _07598_ register_file\[15\]\[9\] _07600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13646__I _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12129_ _06926_ register_file\[3\]\[12\] _06932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08309__A1 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12105__A2 _06912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13302__A1 _07572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07780__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11864__A1 _06770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15055__A1 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15819_ _00207_ clknet_leaf_132_clk register_file\[26\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__A1 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14802__A1 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09340_ _04651_ _04654_ _04655_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11616__A1 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09271_ _04584_ _04587_ _04026_ _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13369__A1 _07708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08222_ _03548_ _03551_ _01101_ _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14030__A2 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11919__A2 _06799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08153_ _03482_ _03483_ _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08796__A1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08084_ _01130_ register_file\[28\]\[27\] _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16024__CLK clknet_leaf_243_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15530__A2 _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12344__A2 _07071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10355__A1 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08986_ _04305_ _04306_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input33_I new_value[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07937_ _02940_ register_file\[12\]\[25\] _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10107__A1 _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13844__A2 _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11855__A1 _06024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10658__A2 register_file\[1\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07868_ _01530_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09607_ _03863_ _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15597__A2 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13291__I _07630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07799_ _03051_ register_file\[1\]\[23\] _03052_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11804__I _06729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09538_ _04582_ register_file\[24\]\[14\] _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09469_ _04576_ register_file\[15\]\[13\] _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12280__A1 _07032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11083__A2 _06269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11500_ _06442_ _06498_ _06540_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12480_ _06990_ _07153_ _07155_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09028__A2 register_file\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11431_ _06373_ _06496_ _06500_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12583__A2 register_file\[22\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14150_ _01411_ register_file\[21\]\[6\] _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13780__A1 _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11362_ _06382_ _06458_ _06459_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_193_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13101_ _07546_ _07544_ _07547_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10313_ _05481_ register_file\[5\]\[25\] _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14081_ _01249_ register_file\[10\]\[5\] _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11293_ _06410_ _06408_ _06411_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15521__A2 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13032_ _07302_ _07494_ _07498_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16517__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10244_ _05531_ _05546_ _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12370__I _07086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10175_ _05471_ _05478_ _05479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10897__A2 _06029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14088__A2 register_file\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14983_ _01649_ _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11846__A1 _06708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13934_ _01451_ _01173_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13865_ _01382_ register_file\[19\]\[3\] _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15604_ _01423_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12816_ _07369_ _07370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_16584_ _00972_ clknet_5_12__leaf_clk register_file\[9\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15691__CLK clknet_leaf_135_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13796_ _01072_ register_file\[26\]\[2\] _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15535_ _03024_ _03033_ _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12271__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11074__A2 _06269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12747_ _07257_ _07322_ _07328_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12678_ _07279_ register_file\[21\]\[19\] _07282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15466_ register_file\[3\]\[21\] _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09019__A2 register_file\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16047__CLK clknet_leaf_245_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14417_ _01921_ _01928_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11629_ _06613_ register_file\[10\]\[17\] _06619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12023__A1 _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15397_ _02895_ _02896_ _02814_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12574__A2 _07208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14348_ _01856_ _01860_ _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14279_ _01790_ _01792_ _01709_ _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15512__A2 register_file\[31\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16197__CLK clknet_leaf_80_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12326__A2 register_file\[25\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13523__A1 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16018_ _00406_ clknet_leaf_229_clk register_file\[6\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10337__A1 _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13376__I _07689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ _04090_ register_file\[6\]\[4\] _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15276__A1 _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14079__A2 _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ _04089_ _04093_ _04094_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10014__B _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15591__I _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_1_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11837__A1 _06698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11624__I _06601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_306_clk_I clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09258__A2 register_file\[30\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09323_ _04622_ _04639_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11065__A2 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _04539_ _04571_ _04298_ net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10812__A2 _06074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14003__A2 _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10684__B _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08205_ _03516_ _03535_ _03303_ _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12014__A1 _06716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09185_ _04497_ _04503_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12565__A2 _07201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13762__A1 _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ _03465_ _03466_ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10576__A1 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08067_ _03068_ register_file\[20\]\[27\] _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12317__A2 register_file\[25\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07992__A2 register_file\[24\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10328__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12190__I _06962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08969_ _03922_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13817__A2 _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11980_ _06682_ _06840_ _06842_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14490__A2 register_file\[18\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10931_ _06069_ _06178_ _06184_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10500__A1 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13650_ _01164_ _01168_ _01170_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10862_ net27 _06133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09249__A2 register_file\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09004__I _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12601_ _07183_ register_file\[22\]\[29\] _07227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12253__A1 _07007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11056__A2 register_file\[28\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13581_ _01088_ _01099_ _01101_ _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ _06076_ _06077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_306_clk clknet_5_1__leaf_clk clknet_leaf_306_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15320_ _02736_ register_file\[30\]\[20\] _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12532_ _07186_ register_file\[22\]\[0\] _07187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10594__B _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12463_ _07137_ _07145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15251_ _02748_ _02752_ _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12005__A1 _06851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14202_ _01623_ _01714_ _01716_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11414_ _06436_ _06486_ _06489_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15182_ _01423_ _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12394_ _07102_ register_file\[24\]\[9\] _07104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09421__A2 register_file\[21\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10567__A1 _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14133_ _01478_ register_file\[30\]\[6\] _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11345_ _06447_ _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15907__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12308__A2 _07050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14064_ _01578_ _01579_ _01494_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11276_ _06398_ _06396_ _06399_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13015_ _07484_ register_file\[17\]\[21\] _07489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11709__I _06081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10227_ _05524_ _05529_ _04026_ _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08932__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10158_ _05460_ _05461_ _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11819__A1 _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10089_ _05386_ _05393_ _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14966_ _02449_ _02470_ _02471_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13917_ _01344_ register_file\[13\]\[3\] _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12492__A1 _07002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14897_ _01038_ _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13848_ _01366_ _01182_ _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14233__A2 register_file\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15430__A1 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12244__A1 _07006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11047__A2 register_file\[28\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16567_ _00955_ clknet_leaf_215_clk register_file\[29\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13779_ _01031_ register_file\[20\]\[2\] _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08753__I _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15518_ _02929_ register_file\[9\]\[22\] _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13992__A1 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_23__f_clk_I clknet_3_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_292_clk_I clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16498_ _00886_ clknet_leaf_175_clk register_file\[15\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12275__I _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15449_ _02939_ _02948_ _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12547__A2 register_file\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10558__A1 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15586__I _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08702__B _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07974__A2 register_file\[16\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09941_ _03919_ _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11619__I _06593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09176__A1 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ _05112_ register_file\[13\]\[19\] _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_230_clk_I clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _04146_ register_file\[6\]\[3\] _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10730__A1 _06024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08754_ _04073_ _04076_ _04078_ _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_245_clk_I clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11286__A2 _06396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08685_ _03975_ _04010_ _03936_ net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_92_clk clknet_5_14__leaf_clk clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__16212__CLK clknet_leaf_157_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11354__I _06449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08151__A2 register_file\[16\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15421__A1 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15270__B _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11038__A2 _06243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09306_ _04556_ register_file\[9\]\[10\] _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09100__A1 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12786__A2 _07350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13983__A1 _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16362__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09651__A2 register_file\[22\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ _04546_ _04554_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13735__A1 _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09168_ _04482_ _04485_ _04486_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10549__A1 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08119_ _03450_ _03374_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11210__A2 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09708__B _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09099_ _04346_ register_file\[6\]\[7\] _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15488__A1 _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11130_ _06130_ _06300_ _06305_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07965__A2 register_file\[1\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14160__A1 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11061_ _06156_ _06257_ _06262_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output64_I net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _05248_ register_file\[23\]\[21\] _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08914__A1 _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13744__I register_file\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14820_ _02316_ _02326_ _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08390__A2 _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14463__A2 register_file\[25\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12474__A1 _07150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14751_ _02258_ register_file\[21\]\[13\] _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11963_ _06665_ _06826_ _06832_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11264__I _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_83_clk clknet_5_11__leaf_clk clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13702_ _01059_ register_file\[25\]\[1\] _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10914_ _06169_ _06174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14682_ _02107_ register_file\[12\]\[12\] _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11894_ _06789_ register_file\[6\]\[14\] _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09890__A2 register_file\[4\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16421_ _00809_ clknet_leaf_73_clk register_file\[17\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12226__A1 _06995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10845_ _06117_ _06118_ _06119_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11029__A2 _06243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07898__B _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13633_ register_file\[7\]\[0\] _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12777__A2 register_file\[20\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16352_ _00740_ clknet_leaf_3_clk register_file\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10776_ _06062_ _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13564_ _01037_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15303_ _02474_ register_file\[24\]\[20\] _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12515_ _07171_ register_file\[23\]\[26\] _07176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16283_ _00671_ clknet_leaf_40_clk register_file\[22\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13495_ _01015_ register_file\[19\]\[0\] _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15234_ _01071_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12446_ _07036_ _07090_ _07133_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12823__I _07361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11201__A2 _06344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15165_ _02667_ register_file\[26\]\[18\] _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12377_ _06967_ _07088_ _07093_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14116_ _01194_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11328_ _06147_ _06436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15096_ _02513_ register_file\[9\]\[17\] _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10960__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11439__I _06497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09158__A1 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11259_ _06386_ _06384_ _06387_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14047_ _01387_ register_file\[28\]\[5\] _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10712__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16235__CLK clknet_leaf_136_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08381__A2 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15998_ _00386_ clknet_leaf_306_clk register_file\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12465__A1 _07142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11268__A2 register_file\[19\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14949_ register_file\[4\]\[15\] _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_74_clk clknet_5_10__leaf_clk clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09330__A1 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08470_ _03775_ _03788_ _03796_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16385__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14206__A2 _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12217__A1 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07892__A1 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09579__I _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12768__A2 register_file\[20\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10779__A1 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09022_ _04059_ register_file\[25\]\[6\] _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14390__A1 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12940__A2 register_file\[18\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09924_ _05229_ _05231_ _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09855_ _04894_ register_file\[24\]\[18\] _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08372__A2 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08806_ _04128_ _04129_ _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09786_ _05092_ _05095_ _04139_ _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11259__A2 _06384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12456__A1 _07138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08737_ _04061_ register_file\[24\]\[2\] _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11084__I _06270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_65_clk clknet_5_10__leaf_clk clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_64_clk_I clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10202__B _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08668_ _03982_ _03993_ _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09872__A2 register_file\[13\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output102_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_199_clk_I clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12908__I _07417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08599_ _03790_ _03814_ _03792_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12759__A2 _07329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10630_ _05925_ _05926_ _05927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_79_clk_I clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10561_ _05668_ register_file\[11\]\[29\] _05859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_122_clk_I clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11431__A2 _06496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12300_ _06969_ _07040_ _07047_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16108__CLK clknet_leaf_193_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13708__A1 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13280_ _07660_ register_file\[14\]\[18\] _07661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10492_ _05527_ register_file\[23\]\[28\] _05791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12231_ _06094_ _06999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09388__A1 _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12643__I _06068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13184__A2 _07601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09438__B _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11195__A1 _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07938__A2 register_file\[13\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12931__A2 _07432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12162_ _06703_ _06950_ _06951_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_137_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10942__A1 _06189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16258__CLK clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _06100_ _06293_ _06295_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14133__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12093_ _06863_ net35 _06909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_17_clk_I clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15921_ _00309_ clknet_leaf_185_clk register_file\[10\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11044_ _06247_ register_file\[28\]\[22\] _06253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12695__A1 _07291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11498__A2 _06534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13474__I _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15852_ _00240_ clknet_leaf_122_clk register_file\[12\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14803_ _02308_ _02309_ _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15783_ _00171_ clknet_leaf_47_clk register_file\[19\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12995_ _07457_ _07477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_56_clk clknet_5_8__leaf_clk clknet_leaf_56_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09312__A1 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12998__A2 register_file\[17\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14734_ _01100_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11946_ _06817_ _06822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09863__A2 register_file\[2\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14665_ _02173_ register_file\[22\]\[12\] _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11877_ _06774_ register_file\[6\]\[7\] _06781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11670__A2 _06641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16404_ _00792_ clknet_leaf_173_clk register_file\[18\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13947__A1 _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13616_ _01131_ _01133_ _01136_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10828_ _06104_ _06096_ _06105_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09615__A2 register_file\[13\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14596_ _02100_ _02105_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16335_ _00723_ clknet_leaf_146_clk register_file\[20\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10338__I _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13547_ _01013_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11422__A2 _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10759_ _06048_ _06049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16266_ _00654_ clknet_leaf_96_clk register_file\[22\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13478_ _00998_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_16_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09379__A1 _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13649__I _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14372__A1 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15217_ _02719_ _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12429_ _07018_ _07119_ _07124_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16197_ _00585_ clknet_leaf_80_clk register_file\[24\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11186__A1 _06082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07929__A2 register_file\[9\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12922__A2 _07432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15148_ _01080_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08051__A1 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10933__A1 _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07970_ _03281_ _03302_ _03303_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_15079_ _02252_ register_file\[18\]\[17\] _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15625__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12686__A1 _07286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09551__A1 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09640_ _04754_ register_file\[29\]\[15\] _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14427__A2 register_file\[10\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10161__A2 register_file\[9\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09571_ _04754_ register_file\[17\]\[14\] _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12438__A1 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_47_clk clknet_5_12__leaf_clk clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08106__A2 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08522_ _03848_ register_file\[18\]\[0\] _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12989__A2 register_file\[17\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11110__A1 _06290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09854__A2 register_file\[25\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13650__A3 _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08453_ _03779_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_180_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08384_ _03711_ _01022_ _01011_ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09606__A2 register_file\[17\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11413__A2 register_file\[26\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08290__A1 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09005_ _04325_ register_file\[21\]\[6\] _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13559__I _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13166__A2 _07584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12463__I _07137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16400__CLK clknet_leaf_160_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11177__A1 _06064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12913__A2 register_file\[18\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10924__A1 _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11079__I _06270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14115__A1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09772__I _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16550__CLK clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09907_ _05213_ _05214_ _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09838_ _05146_ register_file\[29\]\[18\] _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12429__A1 _07018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09769_ _04810_ register_file\[5\]\[17\] _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_38_clk clknet_5_7__leaf_clk clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15091__A2 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11800_ _06734_ register_file\[7\]\[8\] _06735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11101__A1 _06078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12780_ _07347_ register_file\[20\]\[23\] _07348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07856__A1 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11731_ _06687_ register_file\[8\]\[18\] _06688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11652__A2 _06630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13929__A1 _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14450_ _01960_ _01961_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11662_ _06444_ _06594_ _06637_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13401_ _07511_ _07728_ _07733_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10613_ _03868_ register_file\[26\]\[30\] _05910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14381_ _01891_ _01892_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11404__A2 register_file\[26\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12601__A1 _07183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11593_ _06375_ _06592_ _06597_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09947__I _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16120_ _00508_ clknet_leaf_241_clk register_file\[3\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13332_ _07522_ _07690_ _07692_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10544_ _05840_ _05841_ _05842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08281__A1 _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16051_ _00439_ clknet_leaf_231_clk register_file\[5\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16080__CLK clknet_leaf_234_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13157__A2 _07584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__B _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13263_ _07646_ register_file\[14\]\[11\] _07651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10475_ _05640_ register_file\[1\]\[27\] _05775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15002_ _02505_ _02175_ _02506_ _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15648__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12904__A2 register_file\[18\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12214_ _06072_ _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08033__A1 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13194_ _07543_ _07608_ _07609_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10915__A1 _06174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09781__A1 _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12145_ _06686_ _06936_ _06941_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14657__A2 register_file\[18\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12076_ _06899_ net26 _06900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12668__A1 _07267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15798__CLK clknet_leaf_204_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11027_ _06228_ _06243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_110_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09533__A1 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15904_ _00292_ clknet_leaf_7_clk register_file\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15835_ _00223_ clknet_leaf_274_clk register_file\[26\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_29_clk clknet_5_6__leaf_clk clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13093__A1 _07539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15766_ _00154_ clknet_leaf_224_clk register_file\[13\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12978_ _07246_ _07466_ _07467_ _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14717_ _01973_ register_file\[25\]\[13\] _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07847__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11929_ _06767_ register_file\[6\]\[29\] _06811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15697_ _00085_ clknet_leaf_166_clk register_file\[28\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11452__I _06505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14648_ _02149_ _02156_ _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14579_ _01758_ register_file\[23\]\[11\] _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09857__I _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16318_ _00706_ clknet_leaf_30_clk register_file\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14345__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16249_ _00637_ clknet_leaf_193_clk register_file\[23\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11159__A1 _06033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput102 net102 rS[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__14896__A2 register_file\[28\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13699__A3 _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16573__CLK clknet_leaf_304_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08024__A1 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10382__A2 register_file\[13\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12659__A1 _07266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07953_ register_file\[4\]\[25\] _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09524__A1 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13320__A2 register_file\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07884_ _03211_ _03218_ _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09623_ _04669_ register_file\[8\]\[15\] _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14938__I _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15073__A2 register_file\[17\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13084__A1 _07534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09554_ _04667_ register_file\[13\]\[14\] _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08505_ _03831_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12458__I _07137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12831__A1 _07374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09485_ _04797_ _04798_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11634__A2 register_file\[10\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08436_ _03762_ net1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13387__A2 register_file\[29\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08367_ _01182_ register_file\[2\]\[31\] _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_177_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11398__A1 _06419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08298_ _01111_ register_file\[25\]\[30\] _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12193__I _06045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10260_ _03879_ _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_180_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12898__A1 _07246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09763__A1 _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08566__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10191_ _05493_ _05494_ _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15940__CLK clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11570__A1 _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08318__A2 _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13311__A2 _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13950_ _01466_ _01006_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12901_ _07414_ register_file\[18\]\[7\] _07421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11873__A2 register_file\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13881_ _01308_ register_file\[25\]\[3\] _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15620_ _00008_ clknet_leaf_72_clk register_file\[30\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12832_ _07262_ _07377_ _07379_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07829__A1 _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15551_ _02877_ _03047_ _03049_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12368__I _07086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12763_ _07333_ register_file\[20\]\[16\] _07338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11625__A2 register_file\[10\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12822__A1 _07252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16446__CLK clknet_leaf_304_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14502_ _01932_ register_file\[8\]\[10\] _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11714_ _06675_ register_file\[8\]\[13\] _06676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15482_ _02812_ register_file\[18\]\[22\] _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12694_ _06134_ _07293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14575__A1 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14433_ _01603_ register_file\[14\]\[9\] _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13378__A2 _07718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11645_ _06426_ _06623_ _06628_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11389__A1 _06469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08581__I _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14364_ _01876_ _01707_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput15 new_value[13] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08254__A1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16596__CLK clknet_leaf_214_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12050__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput26 new_value[23] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11576_ _06438_ _06582_ _06586_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_183_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13199__I _07582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput37 new_value[4] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10061__A1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16103_ _00491_ clknet_leaf_42_clk register_file\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13315_ _07681_ _07682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10527_ _05563_ register_file\[13\]\[28\] _05826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14295_ _01550_ register_file\[25\]\[8\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16034_ _00422_ clknet_leaf_314_clk register_file\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10458_ _04415_ _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13246_ _07516_ _07632_ _07640_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12889__A1 _07239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09754__A1 _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08557__A2 register_file\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13177_ _07526_ _07594_ _07599_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10389_ _05423_ register_file\[21\]\[26\] _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11561__A1 _06572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08530__B _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12128_ _06670_ _06929_ _06931_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09506__A1 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11447__I _06497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13302__A2 _07670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12059_ _06885_ net18 _06890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11313__A1 _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15055__A2 register_file\[25\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15818_ _00206_ clknet_leaf_104_clk register_file\[26\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13066__A1 _07514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__A2 register_file\[22\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14802__A2 register_file\[25\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15749_ _00137_ clknet_leaf_69_clk register_file\[13\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11616__A2 _06609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12278__I _06155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12813__A1 _07366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09270_ _04585_ _04586_ _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08221_ _03549_ _01094_ _03550_ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14566__A1 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13369__A2 register_file\[29\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09587__I _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08152_ _01111_ register_file\[17\]\[28\] _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12041__A2 _06874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09993__A1 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08083_ _03411_ _03414_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_5_15__f_clk clknet_3_3_0_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09536__B _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11552__A1 _06572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10355__A2 register_file\[24\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16319__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08985_ _04239_ register_file\[28\]\[6\] _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07936_ _03266_ _03269_ _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input26_I new_value[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11855__A2 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07867_ _03199_ _03201_ _02953_ _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13572__I _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16469__CLK clknet_leaf_215_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15046__A2 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09606_ _04917_ register_file\[17\]\[15\] _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08666__I _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09271__B _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07798_ _02877_ _03130_ _03133_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09537_ _04580_ register_file\[25\]\[14\] _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12804__A1 _07362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11092__I _06270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09468_ _04781_ register_file\[14\]\[13\] _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12280__A2 _07024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15499__I _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10291__A1 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14557__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08419_ _03746_ _03657_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09399_ _04711_ _04713_ _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11430_ _06498_ register_file\[12\]\[1\] _06500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08236__A1 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14309__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10043__A1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09984__A1 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11361_ _06454_ register_file\[26\]\[5\] _06459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13100_ _07539_ register_file\[16\]\[16\] _07547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output94_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10312_ _05596_ _05613_ _05614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11292_ _06403_ register_file\[19\]\[16\] _06411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14080_ _01247_ register_file\[11\]\[5\] _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09736__A1 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10243_ _05538_ _05545_ _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13031_ _07455_ register_file\[17\]\[28\] _07498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11543__A1 _06405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10174_ _05474_ _05477_ _04191_ _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11267__I _06068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14982_ _02321_ register_file\[30\]\[16\] _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13933_ _01445_ _01450_ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11846__A2 _06758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13048__A1 _07507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13864_ _01014_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15836__CLK clknet_leaf_279_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15603_ _03099_ _03100_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12815_ _07361_ _07369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12098__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16583_ _00971_ clknet_leaf_49_clk register_file\[9\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13795_ _01313_ register_file\[27\]\[2\] _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15534_ _03029_ _03032_ _02862_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12746_ _07326_ register_file\[20\]\[9\] _07328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12271__A2 _07024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14548__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10282__A1 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15465_ _02964_ register_file\[2\]\[21\] _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_31_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12677_ _06112_ _07281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15986__CLK clknet_leaf_229_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11730__I _06639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14012__A3 _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14416_ _01924_ _01927_ _01671_ _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11628_ _06410_ _06616_ _06618_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15396_ _02812_ register_file\[18\]\[21\] _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12023__A2 _06864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13220__A1 _07570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09200__I _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09975__A1 _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14347_ _01857_ _01858_ _01859_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11559_ _06572_ register_file\[11\]\[21\] _06577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11782__A1 _06722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14278_ _01791_ _01707_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13657__I _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16017_ _00405_ clknet_leaf_229_clk register_file\[6\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13229_ _07583_ register_file\[15\]\[31\] _07629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13523__A2 register_file\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11534__A1 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_260_clk clknet_5_19__leaf_clk clknet_leaf_260_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13287__A1 _07660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08770_ _03876_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13606__B _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11837__A2 _06751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13392__I _07726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09322_ _04629_ _04638_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14539__A1 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12736__I _07321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09253_ _04555_ _04570_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_181_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08204_ _03527_ _03534_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09184_ _04502_ _04294_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12014__A2 _06818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08135_ _03222_ register_file\[25\]\[28\] _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11773__A1 _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16141__CLK clknet_leaf_140_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08066_ _03394_ _03397_ _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_190_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09718__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12471__I _07137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11525__A1 _06550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10328__A2 register_file\[29\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15267__A2 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08941__A2 _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_251_clk clknet_5_16__leaf_clk clknet_leaf_251_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13278__A1 _07548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08968_ _04154_ register_file\[3\]\[5\] _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09780__I _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15859__CLK clknet_leaf_176_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07919_ _03003_ register_file\[20\]\[25\] _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08899_ _03917_ register_file\[2\]\[4\] _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10930_ _06182_ register_file\[2\]\[9\] _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10500__A2 register_file\[7\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10861_ _06130_ _06118_ _06132_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12600_ _07030_ _07222_ _07226_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13580_ _01100_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12253__A2 register_file\[31\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13450__A1 _07560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10792_ net13 _06076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14347__B _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12531_ _07185_ _07186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_40_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12646__I _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15250_ _02749_ _02750_ _02751_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13202__A1 _07612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12462_ _06972_ _07136_ _07144_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10016__A1 _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14201_ _01715_ _01456_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11413_ _06483_ register_file\[26\]\[27\] _06489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15181_ _02682_ _02683_ _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14861__I register_file\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14950__A1 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12393_ _06982_ _07098_ _07103_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11764__A1 _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10567__A2 register_file\[14\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14132_ _01645_ _01475_ _01646_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11344_ _06446_ _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14082__B _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09709__A1 _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14063_ _01405_ register_file\[18\]\[5\] _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11275_ _06391_ register_file\[19\]\[11\] _06399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11516__A1 _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13014_ _07283_ _07487_ _07488_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10226_ _05526_ _05528_ _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_242_clk clknet_5_17__leaf_clk clknet_leaf_242_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10157_ _05192_ register_file\[19\]\[23\] _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08932__A2 register_file\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13269__A1 _07538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10088_ _05389_ _05392_ _04131_ _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14965_ _01194_ _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11819__A2 register_file\[7\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14481__A3 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13916_ _01253_ register_file\[12\]\[3\] _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08696__A1 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12492__A2 _07160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14896_ _02235_ register_file\[28\]\[15\] _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13847_ register_file\[3\]\[2\] _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15430__A2 register_file\[9\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16566_ _00954_ clknet_leaf_215_clk register_file\[29\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12244__A2 _07000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13441__A1 _07550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13778_ _01293_ _01296_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10255__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14257__B _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15517_ _02764_ register_file\[8\]\[22\] _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12556__I _07193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12729_ _07239_ _07312_ _07317_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16497_ _00885_ clknet_leaf_175_clk register_file\[15\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13992__A2 register_file\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16164__CLK clknet_leaf_75_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15194__A1 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15448_ _02943_ _02947_ _02862_ _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09948__A1 _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15379_ _02879_ _02715_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11755__A1 _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10558__A2 register_file\[8\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08620__A1 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15497__A2 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10804__I _06085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09940_ _05117_ register_file\[30\]\[20\] _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12291__I _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09871_ _05145_ _05179_ _04977_ net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_233_clk clknet_5_20__leaf_clk clknet_leaf_233_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_140_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08822_ _04145_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10730__A2 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08753_ _04077_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08684_ _03994_ _04009_ _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08687__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13850__I _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15421__A2 register_file\[30\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14224__A3 _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09305_ _04614_ _04621_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09100__A2 register_file\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10246__A1 _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11994__A1 _06696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09236_ _04549_ _04552_ _04553_ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09167_ _04067_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_33_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08118_ register_file\[5\]\[27\] _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08611__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09098_ _04414_ _04417_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15488__A2 register_file\[22\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08049_ register_file\[3\]\[26\] _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13499__A1 _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15681__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11060_ _06218_ register_file\[28\]\[29\] _06262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14160__A2 register_file\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10011_ _05117_ register_file\[22\]\[21\] _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12171__A1 _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_224_clk clknet_5_21__leaf_clk clknet_leaf_224_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output57_I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16037__CLK clknet_leaf_314_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14750_ _01085_ _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11962_ _06830_ register_file\[5\]\[9\] _06832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08678__A1 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13701_ _01056_ register_file\[24\]\[1\] _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10485__A1 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10913_ _06037_ _06168_ _06173_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14681_ _02186_ _02189_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11893_ _06674_ _06785_ _06790_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16420_ _00808_ clknet_leaf_73_clk register_file\[17\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13632_ _01152_ register_file\[6\]\[0\] _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12226__A2 register_file\[31\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10844_ _06109_ register_file\[30\]\[20\] _06119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13423__A1 _07742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10237__A1 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16351_ _00739_ clknet_leaf_3_clk register_file\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13563_ _01083_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13974__A2 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11280__I _06085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10775_ net41 _06062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15302_ _02763_ _02803_ _02473_ net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11985__A1 _06686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12514_ _07023_ _07174_ _07175_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16282_ _00670_ clknet_leaf_269_clk register_file\[22\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13494_ _01014_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08850__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15233_ _02732_ _02733_ _02734_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14591__I _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12445_ _07087_ register_file\[24\]\[31\] _07133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13726__A2 _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09685__I _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15164_ _01404_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12376_ _07090_ register_file\[24\]\[2\] _07093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14115_ _01622_ _01630_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11327_ _06434_ _06432_ _06435_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15095_ _02349_ register_file\[8\]\[17\] _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13000__I _07465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_305_clk_I clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10960__A2 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14151__A2 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14046_ _01555_ _01561_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11258_ _06378_ register_file\[19\]\[6\] _06387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12162__A1 _06703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_215_clk clknet_5_23__leaf_clk clknet_leaf_215_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10209_ _05506_ _05512_ _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11189_ _06086_ _06337_ _06342_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10712__A2 register_file\[14\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15100__A1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15997_ _00385_ clknet_leaf_307_clk register_file\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14948_ _02451_ _02453_ _02120_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08669__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12465__A2 register_file\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09330__A2 register_file\[27\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14879_ _02385_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12217__A2 _06988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13414__A1 _07524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07892__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16549_ _00937_ clknet_leaf_65_clk register_file\[29\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13965__A2 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09094__A1 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10779__A2 register_file\[30\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15167__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08841__A1 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14715__B _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09021_ _04338_ _04341_ _04201_ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11728__A1 _06684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08713__B _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14390__A2 register_file\[29\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10400__A1 _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09923_ _05230_ register_file\[8\]\[19\] _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12153__A1 _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_206_clk clknet_5_22__leaf_clk clknet_leaf_206_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_86_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09854_ _04892_ register_file\[25\]\[18\] _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11900__A1 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ _04054_ register_file\[27\]\[3\] _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09785_ _05093_ _05094_ _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08736_ _03882_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12456__A2 register_file\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13653__A1 _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09321__A2 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10467__A1 _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08667_ _03985_ _03990_ _03992_ _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07999__B _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13580__I _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13405__A1 _07734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08598_ _03918_ _03921_ _03924_ _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10219__A1 _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12196__I _06049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09085__A1 _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11967__A1 _06830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15158__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08832__A1 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10560_ _05666_ register_file\[10\]\[29\] _05858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09219_ _04533_ _04536_ _04400_ _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13708__A2 register_file\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10491_ _05525_ register_file\[22\]\[28\] _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12230_ _06997_ _06988_ _06998_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09388__A2 register_file\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12392__A1 _07102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11195__A2 register_file\[13\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12161_ _06947_ register_file\[3\]\[25\] _06951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10942__A2 register_file\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11112_ _06290_ register_file\[27\]\[16\] _06295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14133__A2 register_file\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12092_ _03666_ _06866_ _06908_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12144__A1 _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11043_ _06122_ _06250_ _06252_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15920_ _00308_ clknet_leaf_186_clk register_file\[10\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__I _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08899__A1 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_291_clk_I clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15851_ _00239_ clknet_leaf_122_clk register_file\[12\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14802_ _01973_ register_file\[25\]\[14\] _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14436__A3 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15782_ _00170_ clknet_5_14__leaf_clk register_file\[19\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12994_ _07264_ _07473_ _07476_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12447__A2 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14733_ _02239_ _01906_ _02240_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08115__A3 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14586__I _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11945_ _06647_ _06816_ _06821_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13490__I _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14664_ _01089_ _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11876_ _06658_ _06778_ _06780_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16403_ _00791_ clknet_leaf_168_clk register_file\[18\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13615_ _01135_ register_file\[13\]\[0\] _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10827_ _06087_ register_file\[30\]\[17\] _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14595_ _02102_ _02104_ _01859_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11958__A1 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16334_ _00722_ clknet_leaf_145_clk register_file\[20\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15149__A1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13546_ _01064_ _01066_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10758_ net38 _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08823__A1 _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16265_ _00653_ clknet_leaf_96_clk register_file\[22\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13477_ _00997_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_16_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10689_ _03908_ register_file\[19\]\[31\] _05985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15216_ _02717_ _02718_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12428_ _07123_ register_file\[24\]\[23\] _07124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16196_ _00584_ clknet_leaf_76_clk register_file\[24\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11186__A2 _06337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_244_clk_I clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16202__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15147_ _02645_ _02649_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12359_ _07039_ register_file\[25\]\[28\] _07082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10933__A2 register_file\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15321__A1 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14124__A2 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15078_ _02581_ register_file\[19\]\[17\] _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12135__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13665__I _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14029_ _01545_ _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09000__A1 _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_259_clk_I clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12686__A2 _07284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16352__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10697__A1 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09551__A2 register_file\[31\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09570_ _04879_ _04882_ _04118_ _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12438__A2 _07126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08521_ _03847_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11110__A2 register_file\[27\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08452_ _03778_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15388__A1 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08494__I _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08383_ _03705_ _03710_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11949__A1 _06822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10621__A1 _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08290__A2 register_file\[21\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09004_ _03964_ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_178_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15560__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11177__A2 _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12374__A1 _07090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08042__A2 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10924__A2 _06178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15312__A1 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14115__A2 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12126__A1 _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09906_ _05148_ register_file\[28\]\[19\] _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13874__A1 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10688__A1 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09837_ _03840_ _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_19_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12429__A2 _07119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09768_ _05060_ _05077_ _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ _04042_ _04043_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09699_ _05006_ _05009_ _04675_ _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11101__A2 _06286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11823__I _06718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08618__B _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11730_ _06639_ _06687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10860__A1 _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11661_ _06591_ register_file\[10\]\[31\] _06637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14051__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13400_ _07730_ register_file\[9\]\[2\] _07733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10612_ _05907_ _05908_ _05909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14380_ _01550_ register_file\[25\]\[9\] _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08805__A1 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11592_ _06594_ register_file\[10\]\[2\] _06597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13331_ _07686_ register_file\[29\]\[6\] _07692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16225__CLK clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10543_ _03824_ register_file\[28\]\[29\] _05841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08281__A2 register_file\[17\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15030__I register_file\[7\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08353__B _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16050_ _00438_ clknet_leaf_230_clk register_file\[5\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13262_ _07531_ _07649_ _07650_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14354__A2 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15551__A1 _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10474_ _05508_ register_file\[3\]\[27\] _05774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15001_ _02176_ register_file\[23\]\[16\] _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12365__A1 _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12213_ _06985_ _06976_ _06986_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09230__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13193_ _07605_ register_file\[15\]\[15\] _07609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08033__A2 register_file\[6\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10915__A2 register_file\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16375__CLK clknet_leaf_202_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15303__A1 _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12144_ _06940_ register_file\[3\]\[18\] _06941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09781__A2 register_file\[28\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08584__A3 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12117__A1 _06918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13485__I _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12075_ _06862_ _06899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12668__A2 register_file\[21\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13865__A1 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11026_ _06091_ _06236_ _06242_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08336__A3 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15903_ _00291_ clknet_leaf_10_clk register_file\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10679__A1 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15834_ _00222_ clknet_leaf_265_clk register_file\[26\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12977_ _07462_ register_file\[17\]\[5\] _07467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15765_ _00153_ clknet_leaf_217_clk register_file\[13\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11733__I _06112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15205__I register_file\[5\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14716_ _02057_ register_file\[24\]\[13\] _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11928_ _06710_ _06806_ _06810_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15696_ _00084_ clknet_leaf_165_clk register_file\[28\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07847__A2 register_file\[8\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14647_ _02152_ _02155_ _01825_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14042__A1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11859_ _06769_ _06770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_53_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14578_ _01755_ register_file\[22\]\[11\] _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10603__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16317_ _00705_ clknet_leaf_30_clk register_file\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13529_ _01044_ _01046_ _01049_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08272__A2 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_183_clk_I clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16248_ _00636_ clknet_leaf_193_clk register_file\[23\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14345__A2 register_file\[10\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15542__A1 _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12356__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11159__A2 _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_63_clk_I clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput103 net103 rS[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_16179_ _00567_ clknet_5_31__leaf_clk register_file\[25\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07783__A1 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12108__A1 _06649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13395__I _07729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11908__I _06777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08489__I _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07952_ _03283_ _03285_ _02953_ _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12659__A2 _07260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_78_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07883_ _03217_ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_121_clk_I clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ _04667_ register_file\[9\]\[15\] _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15892__CLK clknet_leaf_213_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09553_ _04862_ _04865_ _04183_ _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09288__A1 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13084__A2 _07532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14281__A1 _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15115__I register_file\[7\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11643__I _06590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08504_ _03830_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_64_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11095__A1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09484_ _04663_ register_file\[19\]\[13\] _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07838__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12831__A2 register_file\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_136_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08435_ net2 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_12_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16248__CLK clknet_leaf_193_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14033__A1 _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_16_clk_I clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08366_ _03693_ _01025_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_177_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11398__A2 _06479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12595__A1 _07219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08297_ _01108_ register_file\[24\]\[30\] _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16398__CLK clknet_leaf_144_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08015__A2 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12898__A2 _07418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09763__A2 register_file\[22\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10190_ _05361_ register_file\[15\]\[23\] _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11570__A2 _06582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08399__I register_file\[29\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12900_ _07250_ _07418_ _07420_ _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_189_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13880_ _01056_ register_file\[24\]\[3\] _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12831_ _07374_ register_file\[1\]\[11\] _07379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08348__B _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15550_ _03048_ _02715_ _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11086__A1 _06275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12762_ _07271_ _07336_ _07337_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07829__A2 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12822__A2 _07370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14501_ _01993_ _02011_ _01930_ _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10833__A1 _06109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11713_ _06642_ _06675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15481_ _02646_ register_file\[19\]\[22\] _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14864__I _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12693_ _07290_ _07284_ _07292_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14432_ _01942_ _01775_ _01943_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11644_ _06627_ register_file\[10\]\[23\] _06628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14575__A2 register_file\[20\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15615__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12586__A1 _07016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12384__I _07097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14363_ register_file\[5\]\[8\] _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput16 new_value[14] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08254__A2 register_file\[14\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11575_ _06543_ register_file\[11\]\[28\] _06586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput27 new_value[24] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16102_ _00490_ clknet_leaf_44_clk register_file\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13314_ _07678_ _07681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput38 new_value[5] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10061__A2 register_file\[8\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10526_ _05817_ _05824_ _05825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14294_ _01635_ register_file\[24\]\[8\] _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12338__A1 _07068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16033_ _00421_ clknet_leaf_314_clk register_file\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13245_ _07638_ register_file\[14\]\[4\] _07640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08006__A2 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10457_ _05756_ register_file\[29\]\[27\] _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12889__A2 _07408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09693__I _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13176_ _07598_ register_file\[15\]\[8\] _07599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10388_ _05685_ _05688_ _04045_ _05689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12127_ _06926_ register_file\[3\]\[11\] _06931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12058_ _02455_ _06888_ _06889_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11313__A2 _06420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12510__A1 _07171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11009_ _06060_ _06229_ _06232_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_5_17__f_clk_I clknet_3_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15817_ _00205_ clknet_leaf_105_clk register_file\[26\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14263__A1 _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13066__A2 register_file\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11077__A1 _06271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15748_ _00136_ clknet_leaf_69_clk register_file\[13\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15679_ _00067_ clknet_leaf_19_clk register_file\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08220_ _03320_ register_file\[23\]\[29\] _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16540__CLK clknet_leaf_282_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12577__A1 _07006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08151_ _03243_ register_file\[16\]\[28\] _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09442__A1 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08245__A2 _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09993__A2 register_file\[23\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14318__A2 _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08082_ _03412_ _03413_ _03168_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12329__A1 _07061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14869__A3 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08721__B _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11001__A1 _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14014__I _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08984_ _04237_ register_file\[29\]\[6\] _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13829__A1 _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08012__I _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07935_ _03267_ _03268_ _03108_ _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15554__B _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12501__A1 _07164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07866_ _03200_ _03037_ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08181__A1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09605_ _03860_ _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input19_I new_value[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16070__CLK clknet_leaf_309_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07797_ _03131_ _03132_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11068__A1 _06266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09536_ _04845_ _04848_ _03962_ _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14684__I _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09467_ _03827_ _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_40_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09778__I _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08418_ register_file\[19\]\[31\] _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14557__A2 register_file\[28\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10291__A2 register_file\[23\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ _04712_ register_file\[16\]\[12\] _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15788__CLK clknet_leaf_123_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08349_ _03676_ _03677_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08236__A2 register_file\[30\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10043__A2 register_file\[13\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11240__A1 _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14309__A2 register_file\[30\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11360_ _06457_ _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09984__A2 register_file\[14\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15506__A1 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10311_ _05603_ _05612_ _05613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12932__I _07417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11291_ _06099_ _06410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09727__B _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output87_I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13030_ _07300_ _07494_ _07497_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10242_ _05541_ _05544_ _04873_ _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13532__A3 _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12740__A1 _07250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11543__A2 _06561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10452__I _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10173_ _05475_ _05476_ _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14981_ _02484_ _02318_ _02485_ _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14493__A1 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13932_ _01447_ _01449_ _01273_ _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13863_ _01380_ _01292_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14245__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13048__A2 register_file\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11059__A1 _06152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12814_ _07244_ _07360_ _07368_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15602_ _02929_ register_file\[9\]\[23\] _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16582_ _00970_ clknet_leaf_49_clk register_file\[9\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13794_ _01068_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10806__A1 _06087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14808__B _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12745_ _07254_ _07322_ _07327_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15533_ _03030_ _02945_ _03031_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_5_21__f_clk clknet_3_5_0_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08592__I _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15464_ _01151_ _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12676_ _07278_ _07272_ _07280_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14548__A2 register_file\[24\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12559__A1 _07198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14415_ _01925_ _01757_ _01926_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11627_ _06613_ register_file\[10\]\[16\] _06618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09424__A1 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15395_ _02646_ register_file\[19\]\[21\] _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08227__A2 _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13220__A2 _07622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14346_ _01125_ _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11558_ _06419_ _06575_ _06576_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07986__A1 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11782__A2 register_file\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13938__I _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10509_ _05804_ _05807_ _04191_ _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14277_ register_file\[5\]\[7\] _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11489_ _06531_ register_file\[12\]\[25\] _06535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16016_ _00404_ clknet_leaf_229_clk register_file\[6\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13228_ _07578_ _07586_ _07628_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11534__A2 _06561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12731__A1 _07318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13159_ _07509_ _07584_ _07588_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_170_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14484__A1 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13287__A2 register_file\[14\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13673__I _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08163__A1 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12289__I _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07910__A1 _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09321_ _04635_ _04637_ _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12798__A1 _07308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__A1 _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11470__A1 _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09252_ _04564_ _04569_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10273__A2 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14539__A2 register_file\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08203_ _03533_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09183_ _04498_ _04500_ _04501_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08218__A2 _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09415__A1 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11222__A1 _06148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08134_ _03306_ register_file\[24\]\[28\] _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08007__I _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11773__A2 register_file\[8\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08065_ _03395_ _03396_ _03231_ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07846__I _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16436__CLK clknet_leaf_167_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08967_ _04288_ register_file\[2\]\[5\] _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13278__A2 _07656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13583__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11289__A1 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07918_ _03248_ _03251_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08898_ _04215_ _04218_ _04220_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16586__CLK clknet_leaf_115_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07849_ _03182_ _03183_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10860_ _06131_ register_file\[30\]\[23\] _06132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12789__A1 _07347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09519_ _04832_ register_file\[11\]\[13\] _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12927__I _07406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10791_ _06073_ _06074_ _06075_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13450__A2 _07759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12530_ _07182_ _07185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11461__A1 _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12461_ _07142_ register_file\[23\]\[4\] _07144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14200_ register_file\[3\]\[6\] _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10016__A2 register_file\[16\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11213__A1 _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11412_ _06434_ _06486_ _06488_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15180_ _02513_ register_file\[9\]\[18\] _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12392_ _07102_ register_file\[24\]\[8\] _07103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13758__I _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14131_ _01564_ register_file\[29\]\[6\] _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11764__A2 register_file\[8\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11343_ _06024_ _03794_ _06446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09709__A2 register_file\[13\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14062_ _01313_ register_file\[19\]\[5\] _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11274_ _06077_ _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13013_ _07484_ register_file\[17\]\[20\] _07488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11516__A2 _06544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10225_ _05527_ register_file\[23\]\[24\] _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15258__A3 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10156_ _05190_ register_file\[18\]\[23\] _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13269__A2 _07649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13493__I _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08587__I _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10087_ _05390_ _05391_ _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14964_ _02461_ _02469_ _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13915_ _01428_ _01432_ _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14218__A1 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14895_ _02395_ _02400_ _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09893__A1 _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15953__CLK clknet_leaf_216_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13846_ _01278_ register_file\[2\]\[2\] _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13777_ _01294_ _01295_ _01026_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16565_ _00953_ clknet_leaf_215_clk register_file\[29\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13441__A2 _07752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10989_ _06217_ _06220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15516_ _02991_ _03014_ _02762_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10255__A2 register_file\[26\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12728_ _07314_ register_file\[20\]\[2\] _07317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16496_ _00884_ clknet_leaf_174_clk register_file\[15\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09211__I _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12659_ _07266_ _07260_ _07268_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15447_ _02944_ _02945_ _02946_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09948__A2 register_file\[16\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15378_ register_file\[3\]\[20\] _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11755__A2 register_file\[8\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12952__A1 _07302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14329_ _01841_ register_file\[21\]\[8\] _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08620__A2 register_file\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10092__I _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09870_ _05162_ _05178_ _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08821_ _03777_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08752_ _03815_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08497__I _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14209__A1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08683_ _04003_ _04008_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08687__A2 register_file\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11691__A1 _06658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09636__A1 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09304_ _04617_ _04620_ _04486_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11443__A1 _06502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10246__A2 register_file\[4\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09235_ _03855_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11994__A2 _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15185__A2 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13196__A1 _07546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09166_ _04483_ _04484_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12943__A1 _07293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08117_ _03203_ _03448_ _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09097_ _04416_ register_file\[4\]\[7\] _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08611__A2 register_file\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15826__CLK clknet_leaf_169_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08048_ _03380_ register_file\[2\]\[26\] _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10010_ _05314_ _05315_ _05316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12171__A2 register_file\[3\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09999_ _03776_ _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10182__A1 _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15976__CLK clknet_leaf_297_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14999__A2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13120__A1 _07551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11961_ _06662_ _06826_ _06831_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09875__A1 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10912_ _06170_ register_file\[2\]\[2\] _06173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13700_ _01211_ _01219_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14680_ _02187_ _02188_ _01859_ _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11682__A1 _06650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10485__A2 register_file\[19\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11892_ _06789_ register_file\[6\]\[13\] _06790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13631_ _01151_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12657__I _07234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10843_ _06051_ _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_77_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13423__A2 register_file\[9\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13562_ _01034_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16350_ _00738_ clknet_leaf_303_clk register_file\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10774_ _06060_ _06052_ _06061_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15301_ _02781_ _02802_ _02471_ _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12513_ _07171_ register_file\[23\]\[25\] _07175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11985__A2 _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16281_ _00669_ clknet_leaf_193_clk register_file\[22\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10177__I _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13493_ _01013_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_160_clk clknet_5_31__leaf_clk clknet_leaf_160_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__A2 register_file\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16601__CLK clknet_leaf_257_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09966__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15232_ _02403_ register_file\[21\]\[19\] _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12444_ _07034_ _07090_ _07132_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15189__B _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13488__I _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12934__A1 _07283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15163_ _02581_ register_file\[27\]\[18\] _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09187__B _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12375_ _06965_ _07088_ _07092_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10905__I _06167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14114_ _01629_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11326_ _06427_ register_file\[19\]\[26\] _06435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15094_ _02574_ _02597_ _02347_ _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14687__A1 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10126__B _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14045_ _01556_ _01558_ _01560_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11257_ _06055_ _06386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10208_ _05511_ _05309_ _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12162__A2 _06950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11188_ _06341_ register_file\[13\]\[13\] _06342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11736__I _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10139_ _05443_ _05309_ _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15996_ _00384_ clknet_5_4__leaf_clk register_file\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13111__A1 _07553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14947_ _02452_ _02203_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09866__A1 _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08669__A2 register_file\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13951__I _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13662__A2 _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11673__A1 _06645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16131__CLK clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14878_ _02383_ _02384_ _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09618__A1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13829_ _01143_ register_file\[15\]\[2\] _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11471__I _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13414__A2 _07738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16548_ _00936_ clknet_leaf_69_clk register_file\[29\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09094__A2 register_file\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16281__CLK clknet_leaf_193_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_151_clk clknet_5_30__leaf_clk clknet_leaf_151_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16479_ _00867_ clknet_leaf_6_clk register_file\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08841__A2 register_file\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13178__A1 _07598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ _04339_ _04340_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15849__CLK clknet_leaf_111_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12925__A1 _07429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11728__A2 _06680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10815__I _06094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10400__A2 register_file\[8\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14678__A1 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15999__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09922_ _03882_ _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13350__A1 _07701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12153__A2 register_file\[3\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09853_ _05154_ _05161_ _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10164__A1 _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11900__A2 _06792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ _04052_ register_file\[26\]\[3\] _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09784_ _05025_ register_file\[31\]\[17\] _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08735_ _04059_ register_file\[25\]\[2\] _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13653__A2 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08666_ _03991_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10467__A2 register_file\[24\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11664__A1 _06216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16096__D _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08597_ _03923_ register_file\[1\]\[0\] _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13405__A2 register_file\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08176__B _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11416__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09085__A2 register_file\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11967__A2 register_file\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_142_clk clknet_5_27__leaf_clk clknet_leaf_142_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__15158__A2 register_file\[24\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13169__A1 _07590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09218_ _04534_ _04535_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10490_ _05787_ _05788_ _05789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12916__A1 _07429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09149_ _04464_ _04467_ _04400_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12392__A2 register_file\[24\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12160_ _06921_ _06950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_194_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11111_ _06095_ _06293_ _06294_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16004__CLK clknet_leaf_314_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09735__B _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12091_ _06863_ net34 _06908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15330__A2 _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08348__A1 _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13341__A1 _07694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11042_ _06247_ register_file\[28\]\[21\] _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11556__I _06553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08899__A2 register_file\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15850_ _00238_ clknet_leaf_111_clk register_file\[12\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16154__CLK clknet_leaf_269_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14801_ _02057_ register_file\[24\]\[14\] _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15781_ _00169_ clknet_leaf_66_clk register_file\[19\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12993_ _07470_ register_file\[17\]\[12\] _07476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14732_ _02071_ register_file\[31\]\[13\] _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11655__A1 _06591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11944_ _06818_ register_file\[5\]\[2\] _06821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14663_ _02170_ _01840_ _02171_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11875_ _06774_ register_file\[6\]\[6\] _06780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11291__I _06099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16402_ _00790_ clknet_leaf_159_clk register_file\[18\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10826_ _06103_ _06104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11407__A1 _06429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13614_ _01134_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14594_ _02103_ register_file\[10\]\[11\] _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16333_ _00721_ clknet_leaf_142_clk register_file\[20\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15149__A2 register_file\[20\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13545_ _01065_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10757_ _06046_ _06027_ _06047_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08823__A2 register_file\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16264_ _00652_ clknet_leaf_91_clk register_file\[22\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13476_ net6 _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_173_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10688_ _03905_ register_file\[18\]\[31\] _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12907__A1 _07257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12427_ _07086_ _07123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15215_ _02634_ register_file\[1\]\[18\] _02635_ _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14107__I _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16195_ _00583_ clknet_leaf_71_clk register_file\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15146_ _02647_ _02648_ _02399_ _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12358_ _07028_ _07078_ _07081_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11309_ _06415_ register_file\[19\]\[21\] _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15077_ _01119_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15321__A2 register_file\[31\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12289_ _07039_ _07040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12135__A2 _06929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13332__A1 _07522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14028_ _01543_ _01544_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10146__A1 _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13883__A2 _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11894__A1 _06789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15979_ _00367_ clknet_leaf_250_clk register_file\[7\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14832__A1 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08520_ _03806_ _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11646__A1 _06627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08451_ _03777_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_64_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13399__A1 _07509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08382_ _03707_ _03709_ _01159_ _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15671__CLK clknet_leaf_224_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14060__A2 _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12071__A1 _06892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_124_clk clknet_5_24__leaf_clk clknet_leaf_124_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09003_ _04315_ _04322_ _04323_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16027__CLK clknet_leaf_252_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15560__A2 register_file\[24\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12374__A2 register_file\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10385__A1 _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12760__I _07321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12126__A2 _06929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13323__A1 _07686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09905_ _05146_ register_file\[29\]\[19\] _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10137__A1 _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13874__A2 register_file\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09836_ _05129_ _05144_ _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11885__A1 _06782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10688__A2 register_file\[18\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08750__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09767_ _05069_ _05076_ _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11637__A1 _06620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08718_ _03851_ register_file\[15\]\[2\] _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09698_ _05007_ _05008_ _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_2__f_clk clknet_3_0_0_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08502__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08649_ _03952_ _03974_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15379__A2 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_304_clk_I clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12000__I _06825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11660_ _06442_ _06594_ _06636_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10860__A2 register_file\[30\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14051__A2 register_file\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10611_ _03864_ register_file\[24\]\[30\] _05908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_115_clk clknet_5_13__leaf_clk clknet_leaf_115_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11591_ _06373_ _06592_ _06596_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08805__A2 register_file\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15311__I _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13330_ _07518_ _07690_ _07691_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10542_ _03821_ register_file\[29\]\[29\] _05840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15000__A1 _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13261_ _07646_ register_file\[14\]\[10\] _07650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10473_ _05637_ register_file\[2\]\[27\] _05773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12212_ _06983_ register_file\[31\]\[9\] _06986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15000_ _02173_ register_file\[22\]\[16\] _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12365__A2 register_file\[25\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13192_ _07593_ _07608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_68_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09230__A2 register_file\[16\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10376__A1 _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12670__I _06103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12143_ _06910_ _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15303__A2 register_file\[24\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12117__A2 register_file\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12074_ _03040_ _06895_ _06898_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10128__A1 _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13865__A2 register_file\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11025_ _06240_ register_file\[28\]\[14\] _06242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15902_ _00290_ clknet_leaf_303_clk register_file\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11876__A1 _06658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15067__A1 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15833_ _00221_ clknet_leaf_263_clk register_file\[26\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14597__I _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11628__A1 _06410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08595__I _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15764_ _00152_ clknet_leaf_177_clk register_file\[13\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12976_ _07465_ _07466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15694__CLK clknet_leaf_152_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14715_ _02181_ _02223_ _02056_ net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11927_ _06767_ register_file\[6\]\[28\] _06810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15695_ _00083_ clknet_leaf_152_clk register_file\[28\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14646_ _02153_ _01906_ _02154_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11858_ _06766_ _06769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_18_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14546__B _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10809_ _06089_ _06090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12053__A1 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14577_ _02085_ _01840_ _02086_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11789_ _06726_ register_file\[7\]\[4\] _06728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16316_ _00704_ clknet_leaf_278_clk register_file\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11800__A1 _06734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10603__A2 register_file\[9\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13528_ _01048_ register_file\[23\]\[0\] _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16247_ _00635_ clknet_leaf_190_clk register_file\[23\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10365__I _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13459_ _07763_ register_file\[9\]\[26\] _07768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12356__A2 _07078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput104 net104 rS[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_16178_ _00566_ clknet_leaf_155_clk register_file\[25\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12580__I _07193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15129_ _02462_ _02630_ _02632_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13305__A1 _07631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12108__A2 _06912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07783__A2 register_file\[6\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08980__A1 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07951_ _03284_ _03037_ _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10119__A1 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07882_ _03215_ _03216_ _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09621_ _04929_ _04932_ _03877_ _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09552_ _04863_ _04864_ _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14300__I _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08503_ _03783_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_70_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11095__A2 register_file\[27\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ _04661_ register_file\[18\]\[13\] _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12292__A1 _07042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08434_ _03721_ _03761_ net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15230__A1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14033__A2 register_file\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12755__I _07313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08365_ _00995_ register_file\[3\]\[31\] _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14584__A3 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15131__I _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08799__A1 _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08296_ _03617_ _03624_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09460__A2 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14336__A3 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15533__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10358__A1 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13586__I _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15297__A1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08723__A1 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09819_ _05124_ _05127_ _04655_ _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10530__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12830_ _07259_ _07377_ _07378_ _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_243_clk_I clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12761_ _07333_ register_file\[20\]\[15\] _07337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11086__A2 register_file\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12283__A1 _07034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14500_ _02003_ _02010_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11712_ _06085_ _06674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15480_ _02977_ _02978_ _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12692_ _07291_ register_file\[21\]\[23\] _07292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15221__A1 _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14431_ _01776_ register_file\[13\]\[9\] _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12035__A1 _06870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11643_ _06590_ _06627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12586__A2 _07215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13783__A1 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14362_ _01531_ _01874_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11574_ _06436_ _06582_ _06585_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10597__A1 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 new_value[15] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16101_ _00489_ clknet_leaf_54_clk register_file\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput28 new_value[25] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10525_ _05820_ _05823_ _03816_ _05824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput39 new_value[6] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13313_ _07679_ _07680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14293_ _01763_ _01806_ _01634_ net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_156_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12338__A2 register_file\[25\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16032_ _00420_ clknet_leaf_1_clk register_file\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13244_ _07513_ _07632_ _07639_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_170_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10456_ _03765_ _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13496__I _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13175_ _07585_ _07598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16492__CLK clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10387_ _05686_ _05687_ _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12126_ _06667_ _06929_ _06930_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08962__A1 _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10134__B _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11849__A1 _06719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12057_ _06885_ net17 _06889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08714__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12510__A2 register_file\[23\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11008_ _06225_ register_file\[28\]\[7\] _06232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14120__I _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15816_ _00204_ clknet_leaf_107_clk register_file\[26\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14263__A2 register_file\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15747_ _00135_ clknet_leaf_54_clk register_file\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12274__A1 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12959_ _06316_ _03854_ _07454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15678_ _00066_ clknet_leaf_24_clk register_file\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12575__I _07182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14629_ _02130_ _02138_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08274__B _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12577__A2 _07208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08150_ _03473_ _03480_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09442__A2 register_file\[24\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10588__A1 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08081_ _03084_ register_file\[26\]\[27\] _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15515__A2 _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09884__I _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12329__A2 register_file\[25\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11001__A2 _06219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15279__A1 _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ _04300_ _04303_ _03962_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13829__A2 register_file\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07934_ _02936_ register_file\[10\]\[25\] _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08705__A1 _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12501__A2 register_file\[23\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07865_ register_file\[7\]\[24\] _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10512__A1 _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16215__CLK clknet_leaf_197_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09604_ _04911_ _04915_ _03796_ _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07796_ _01155_ _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14254__A2 _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11068__A2 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09535_ _04846_ _04847_ _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14965__I _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__A1 _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09466_ _04778_ _04779_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14006__A2 _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08417_ _03706_ register_file\[18\]\[31\] _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09397_ _03772_ _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08348_ _03459_ register_file\[1\]\[30\] _01198_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15506__A2 register_file\[29\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _03571_ _03608_ _03305_ net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10310_ _05606_ _05611_ _04873_ _05612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_193_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07995__A2 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11290_ _06407_ _06408_ _06409_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10241_ _05542_ _05543_ _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14190__A1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10733__I _06025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08944__A1 _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12740__A2 _07322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10172_ _05275_ register_file\[27\]\[23\] _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10751__A1 _06042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14980_ _02403_ register_file\[29\]\[16\] _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14493__A2 register_file\[20\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13931_ _01448_ _01271_ _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10503__A1 _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08172__A2 _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_9__f_clk_I clknet_3_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_182_clk_I clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13862_ _01379_ _01006_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15442__A1 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15601_ _02764_ register_file\[8\]\[23\] _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12256__A1 _07007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11059__A2 _06257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12813_ _07366_ register_file\[1\]\[4\] _07368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16581_ _00969_ clknet_leaf_57_clk register_file\[9\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_309_clk clknet_5_1__leaf_clk clknet_leaf_309_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_34_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_62_clk_I clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13793_ _01311_ _01225_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15532_ _02859_ register_file\[15\]\[22\] _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12744_ _07326_ register_file\[20\]\[8\] _07327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10806__A2 register_file\[30\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_197_clk_I clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12008__A1 _06710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15463_ _02962_ _02793_ _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12675_ _07279_ register_file\[21\]\[18\] _07280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15732__CLK clknet_leaf_177_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12559__A2 register_file\[22\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14414_ _01758_ register_file\[23\]\[9\] _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13756__A1 _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11626_ _06407_ _06616_ _06617_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15394_ _02893_ _01292_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09424__A2 register_file\[22\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14345_ _01684_ register_file\[10\]\[8\] _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09918__B _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11557_ _06572_ register_file\[11\]\[20\] _06576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10508_ _05805_ _05806_ _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11488_ _06505_ _06534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15882__CLK clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14276_ _01531_ _01789_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09188__A1 _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16015_ _00403_ clknet_leaf_244_clk register_file\[6\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13227_ _07583_ register_file\[15\]\[30\] _07628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10439_ _05674_ register_file\[12\]\[27\] _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_135_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12731__A2 register_file\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13158_ _07586_ register_file\[15\]\[1\] _07588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16238__CLK clknet_leaf_145_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12109_ _06918_ register_file\[3\]\[4\] _06920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13089_ _07506_ _07539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_15_clk_I clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08163__A2 register_file\[22\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16388__CLK clknet_leaf_75_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07910__A2 register_file\[16\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12247__A1 _07009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14787__A3 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09320_ _04636_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09112__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12798__A2 _07314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__A2 _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09251_ _04568_ _04294_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11470__A2 _06520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08202_ _03531_ _03532_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09182_ _04291_ register_file\[1\]\[8\] _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08133_ _03425_ _03464_ _03305_ net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11222__A2 _06358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07977__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08064_ _03229_ register_file\[18\]\[27\] _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10981__A1 _06167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09179__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14172__A1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08926__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08023__I _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13864__I _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08966_ _03916_ _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_4706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input31_I new_value[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12486__A1 _07157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07917_ _03249_ _03250_ _03168_ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11384__I _06457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10502__B _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08897_ _04219_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_95_clk clknet_5_15__leaf_clk clknet_leaf_95_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08154__A2 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07848_ _02929_ register_file\[9\]\[24\] _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15755__CLK clknet_leaf_136_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07779_ _02859_ register_file\[15\]\[23\] _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08693__I _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09518_ _04148_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10790_ _06065_ register_file\[30\]\[10\] _06075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11461__A2 _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09449_ _04556_ register_file\[13\]\[12\] _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12460_ _06969_ _07136_ _07143_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11411_ _06483_ register_file\[26\]\[26\] _06488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12410__A1 _06999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12391_ _07089_ _07102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11213__A2 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14130_ _01387_ register_file\[28\]\[6\] _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11342_ _06444_ _06371_ _06445_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10972__A1 _06144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11273_ _06395_ _06396_ _06397_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14061_ _01576_ _01490_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13012_ _07465_ _07487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10224_ _03870_ _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09590__A1 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10155_ _05457_ _05458_ _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08868__I _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14466__A2 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16530__CLK clknet_leaf_175_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12477__A1 _07150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10086_ _05192_ register_file\[27\]\[22\] _05391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14963_ _02468_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11294__I _06103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_86_clk clknet_5_11__leaf_clk clknet_leaf_86_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09342__A1 _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08145__A2 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13914_ _01429_ _01430_ _01431_ _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14894_ _02396_ _02398_ _02399_ _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15415__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14218__A2 register_file\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12229__A1 _06995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13845_ _01363_ _01173_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16564_ _00952_ clknet_leaf_210_clk register_file\[29\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13776_ _01019_ register_file\[18\]\[2\] _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10988_ _06218_ _06219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_128_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15515_ _03002_ _03013_ _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12727_ _07237_ _07312_ _07316_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16495_ _00883_ clknet_leaf_188_clk register_file\[15\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15446_ _02859_ register_file\[15\]\[21\] _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12658_ _07267_ register_file\[21\]\[13\] _07268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12401__A1 _07102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11609_ _06390_ _06602_ _06607_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15377_ _02548_ register_file\[2\]\[20\] _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_8_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12589_ _07018_ _07215_ _07220_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_10_clk clknet_5_3__leaf_clk clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07959__A2 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14328_ _01085_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12952__A2 _07446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08081__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16060__CLK clknet_leaf_293_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10373__I _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14259_ _01688_ register_file\[12\]\[7\] _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15628__CLK clknet_leaf_135_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08908__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08384__A2 _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08820_ _04142_ _04143_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08778__I _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12468__A1 _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08751_ _04074_ _04075_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_77_clk clknet_5_10__leaf_clk clknet_leaf_77_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_113_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15778__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09333__A1 _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08682_ _04007_ _03929_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14209__A2 register_file\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11140__A1 _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11691__A2 _06656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13968__A1 _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09303_ _04618_ _04619_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09234_ _04550_ _04551_ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14393__A1 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09165_ _04348_ register_file\[27\]\[8\] _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13196__A2 _07608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08116_ register_file\[4\]\[27\] _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12943__A2 _07439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09096_ _04415_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10954__A1 _06196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11379__I _06449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14145__A1 _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08047_ _01151_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16553__CLK clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13594__I _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09572__A1 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09998_ _05173_ register_file\[3\]\[20\] _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10182__A2 register_file\[6\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12459__A1 _07142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08949_ _04269_ _04270_ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_68_clk clknet_5_10__leaf_clk clknet_leaf_68_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11960_ _06830_ register_file\[5\]\[8\] _06831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11131__A1 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14639__B _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10911_ _06033_ _06168_ _06172_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07886__A1 _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11891_ _06769_ _06789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11682__A2 register_file\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08637__B _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13630_ _01014_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13959__A1 _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10842_ _06116_ _06117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14620__A2 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12631__A1 _07242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10458__I _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13561_ _01081_ register_file\[28\]\[0\] _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10773_ _06042_ register_file\[30\]\[7\] _06061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15300_ _02794_ _02801_ _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12512_ _07145_ _07174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_73_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16280_ _00668_ clknet_leaf_191_clk register_file\[22\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13492_ _00997_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15176__A3 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15231_ _01083_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14384__A1 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16083__CLK clknet_leaf_231_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12673__I _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12443_ _07087_ register_file\[24\]\[30\] _07132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11198__A1 _06104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14923__A3 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12934__A2 _07439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15162_ _02664_ _01225_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08063__A1 _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12374_ _07090_ register_file\[24\]\[1\] _07092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10945__A1 _06189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14113_ _01627_ _01628_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14136__A1 _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07810__A1 _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11325_ _06143_ _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15093_ _02585_ _02596_ _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14044_ _01559_ _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11256_ _06382_ _06384_ _06385_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08366__A2 _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10207_ _05507_ _05509_ _05510_ _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_45_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11187_ _06321_ _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15920__CLK clknet_leaf_186_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11370__A1 _06462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10138_ _05440_ _05441_ _05442_ _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10142__B _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15995_ _00383_ clknet_leaf_288_clk register_file\[7\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_59_clk clknet_5_8__leaf_clk clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09315__A1 _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13111__A2 _07544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10069_ _05306_ register_file\[1\]\[21\] _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14946_ register_file\[7\]\[15\] _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11122__A1 _06297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09866__A2 register_file\[1\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07877__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14877_ _02217_ register_file\[1\]\[14\] _02218_ _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11673__A2 _06641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12870__A1 _07300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13828_ _01139_ register_file\[14\]\[2\] _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09618__A2 register_file\[14\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16547_ _00935_ clknet_leaf_18_clk register_file\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13759_ _01278_ register_file\[2\]\[1\] _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__16426__CLK clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16478_ _00866_ clknet_leaf_305_clk register_file\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13679__I _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15429_ _01013_ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09378__B _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11189__A1 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12925__A2 register_file\[18\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16576__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10936__A1 _06078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11199__I _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14127__A1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09921_ _05228_ register_file\[9\]\[19\] _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12689__A1 _07288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09554__A1 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10831__I _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13350__A2 register_file\[29\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09852_ _05157_ _05160_ _04017_ _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11361__A1 _06454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08803_ _04123_ _04126_ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09783_ _05023_ register_file\[30\]\[17\] _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09306__A1 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08109__A2 _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08734_ _03879_ _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11113__A1 _06100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08665_ _03836_ _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12861__A1 _07290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11664__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08596_ _03922_ _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11416__A2 _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12613__A1 _07235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08293__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09217_ _04259_ register_file\[23\]\[9\] _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13169__A2 register_file\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09288__B _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12916__A2 register_file\[18\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09148_ _04465_ _04466_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10227__B _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09079_ _04397_ _04398_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11110_ _06290_ register_file\[27\]\[15\] _06294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14669__A2 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12090_ _03593_ _06902_ _06907_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11041_ _06117_ _06250_ _06251_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09545__A1 _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08348__A2 register_file\[1\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13341__A2 register_file\[29\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output62_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11352__A1 _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14800_ _02266_ _02307_ _02056_ net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15780_ _00168_ clknet_leaf_66_clk register_file\[19\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12992_ _07262_ _07473_ _07475_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14731_ _01904_ register_file\[30\]\[13\] _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07859__A1 _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11943_ _06645_ _06816_ _06820_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16449__CLK clknet_leaf_54_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14662_ _01841_ register_file\[21\]\[12\] _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11874_ _06654_ _06778_ _06779_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16401_ _00789_ clknet_leaf_160_clk register_file\[18\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13613_ _01037_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11407__A2 _06479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10825_ _06102_ _06103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12604__A1 _07034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14593_ _01122_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_186_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16332_ _00720_ clknet_leaf_141_clk register_file\[20\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13544_ net9 _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10756_ _06042_ register_file\[30\]\[4\] _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10091__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14357__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16263_ _00651_ clknet_leaf_91_clk register_file\[22\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13475_ _00995_ register_file\[16\]\[0\] _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10687_ _05981_ _05982_ _05983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15214_ _02462_ _02713_ _02716_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12426_ _07016_ _07119_ _07122_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12907__A2 _07418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16194_ _00582_ clknet_leaf_70_clk register_file\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10918__A1 _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09784__A1 _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15145_ _02397_ register_file\[18\]\[18\] _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12357_ _07075_ register_file\[25\]\[27\] _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11591__A1 _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11308_ _06121_ _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15076_ _02579_ _02249_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12288_ _07038_ _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11747__I _06639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13332__A2 _07690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14027_ _01369_ register_file\[1\]\[4\] _01371_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11239_ _06032_ _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10146__A2 register_file\[28\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11343__A1 _06024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15609__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15085__A2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15978_ _00366_ clknet_leaf_291_clk register_file\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07960__I _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14832__A2 register_file\[20\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14929_ _02101_ register_file\[11\]\[15\] _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12843__A1 _07381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08450_ _03776_ net1 _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15816__CLK clknet_leaf_107_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13399__A2 _07728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08381_ _03708_ _03657_ _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10082__A1 _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10826__I _06103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15966__CLK clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14899__A2 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09002_ _04017_ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_178_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08027__A1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13020__A1 _07491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10909__A1 _06021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09775__A1 _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10385__A2 register_file\[14\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11582__A1 _06444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09904_ _05196_ _05211_ _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13323__A2 register_file\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10137__A2 register_file\[1\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09835_ _05136_ _05143_ _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15076__A2 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09766_ _05072_ _05075_ _04900_ _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13087__A1 _07536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08966__I _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08717_ _03848_ register_file\[14\]\[2\] _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12834__A1 _07264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12488__I _07145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09697_ _04939_ register_file\[31\]\[16\] _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08502__A2 register_file\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08648_ _03963_ _03973_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14587__A1 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output100_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13821__B _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08579_ _03905_ register_file\[6\]\[0\] _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10610_ _03861_ register_file\[25\]\[30\] _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12062__A2 _06888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11590_ _06594_ register_file\[10\]\[1\] _06596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10073__A1 _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10541_ _05810_ _05839_ _05647_ net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13112__I _06115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15000__A2 register_file\[22\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08018__A1 _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13011__A1 _07281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13260_ _07641_ _07649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_148_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10472_ _05768_ _05771_ _04068_ _05772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12211_ _06068_ _06985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13191_ _07541_ _07601_ _07607_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11573__A1 _06579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10376__A2 register_file\[30\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16121__CLK clknet_leaf_241_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12142_ _06684_ _06936_ _06939_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15039__I _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14511__A1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12073_ _06892_ net25 _06898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10128__A2 register_file\[9\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11024_ _06086_ _06236_ _06241_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15901_ _00289_ clknet_leaf_280_clk register_file\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15483__B _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11876__A2 _06778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15067__A2 register_file\[31\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15832_ _00220_ clknet_leaf_260_clk register_file\[26\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15839__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15763_ _00151_ clknet_leaf_177_clk register_file\[13\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12825__A1 _07254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12975_ _07457_ _07465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11628__A2 _06616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10420__B _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14714_ _02200_ _02222_ _02054_ _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11926_ _06708_ _06806_ _06809_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15694_ _00082_ clknet_leaf_152_clk register_file\[28\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14578__A1 _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14645_ _02071_ register_file\[31\]\[12\] _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13731__B _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11857_ _06767_ _06768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15989__CLK clknet_leaf_233_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10808_ net16 _06089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14576_ _01841_ register_file\[21\]\[11\] _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13250__A1 _07518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12053__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11788_ _06649_ _06720_ _06727_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10064__A1 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16315_ _00703_ clknet_leaf_272_clk register_file\[21\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13527_ _01047_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_158_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14118__I _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10739_ _06032_ _06033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11800__A2 register_file\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16246_ _00634_ clknet_leaf_183_clk register_file\[23\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13002__A1 _07271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13458_ _07567_ _07766_ _07767_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09757__A1 _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12409_ _07109_ register_file\[24\]\[15\] _07113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16177_ _00565_ clknet_leaf_155_clk register_file\[25\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput105 net105 rS[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_13389_ _07679_ register_file\[29\]\[31\] _07725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11564__A1 _06579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15128_ _02631_ _02300_ _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12082__B _06903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09509__A1 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14502__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13305__A2 register_file\[14\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15059_ _02230_ register_file\[27\]\[17\] _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07950_ register_file\[7\]\[25\] _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08980__A2 register_file\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11316__A1 _06427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10119__A2 register_file\[13\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11867__A2 register_file\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07881_ _03051_ register_file\[1\]\[24\] _03052_ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15058__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09620_ _04930_ _04931_ _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13069__A1 _07514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14805__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09551_ _04663_ register_file\[31\]\[14\] _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08502_ _03828_ register_file\[22\]\[0\] _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09482_ _04794_ _04795_ _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08433_ _03760_ _01105_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15412__I _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15230__A2 register_file\[20\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08248__A1 _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13241__A1 _07511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08364_ _03691_ _01394_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08799__A2 register_file\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13792__A2 _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08295_ _03620_ _03623_ _01101_ _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16144__CLK clknet_leaf_156_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15568__B _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14472__B _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11555__A1 _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10358__A2 register_file\[27\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08470__B _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07865__I register_file\[7\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16294__CLK clknet_leaf_80_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15297__A2 register_file\[1\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_281_clk clknet_5_4__leaf_clk clknet_leaf_281_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11307__A1 _06419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09818_ _05125_ _05126_ _05127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08723__A2 _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09749_ _05055_ _05058_ _04382_ _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12807__A1 _07237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12760_ _07321_ _07336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12283__A2 _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13480__A1 _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11711_ _06672_ _06668_ _06673_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12691_ _07231_ _07291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14430_ _01688_ register_file\[12\]\[9\] _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11642_ _06424_ _06623_ _06626_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12035__A2 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09320__I _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10046__A1 _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14980__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14361_ register_file\[4\]\[8\] _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13783__A2 register_file\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11573_ _06579_ register_file\[11\]\[27\] _06585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16100_ _00488_ clknet_leaf_54_clk register_file\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11794__A1 _06654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput18 new_value[16] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13312_ _07678_ _07679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10524_ _05821_ _05822_ _05823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 new_value[26] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14292_ _01783_ _01805_ _01632_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09739__A1 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16031_ _00419_ clknet_leaf_0_clk register_file\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12681__I _07247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14732__A1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13243_ _07638_ register_file\[14\]\[3\] _07639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10455_ _05749_ _05754_ _05421_ _05755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_182_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11546__A1 _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13174_ _07524_ _07594_ _07597_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08411__A1 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10386_ _05418_ register_file\[15\]\[26\] _05687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11297__I _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15288__A2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12125_ _06926_ register_file\[3\]\[10\] _06930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08962__A2 register_file\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_272_clk clknet_5_7__leaf_clk clknet_leaf_272_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13299__A1 _07667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15661__CLK clknet_leaf_142_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13838__A3 _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12056_ _06873_ _06888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11849__A2 register_file\[7\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11007_ _06056_ _06229_ _06231_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15815_ _00203_ clknet_leaf_107_clk register_file\[26\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16017__CLK clknet_leaf_229_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15746_ _00134_ clknet_leaf_53_clk register_file\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12274__A2 _07024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12958_ _07308_ _07410_ _07453_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11909_ _06796_ register_file\[6\]\[20\] _06800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15677_ _00065_ clknet_leaf_32_clk register_file\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11760__I _06147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12889_ _07239_ _07408_ _07413_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16167__CLK clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14628_ _02137_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13223__A1 _07583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10037__A1 _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09978__A1 _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14971__A1 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14559_ _02067_ _01901_ _02068_ _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13774__A2 _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_26__f_clk_I clknet_3_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11785__A1 _06647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10588__A2 register_file\[5\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08080_ _01120_ register_file\[27\]\[27\] _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08650__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15388__B _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16229_ _00617_ clknet_leaf_78_clk register_file\[23\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14723__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09386__B _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11537__A1 _06558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_263_clk clknet_5_18__leaf_clk clknet_leaf_263_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08982_ _04301_ _04302_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_303_clk_I clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07933_ _02934_ register_file\[11\]\[25\] _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08705__A2 register_file\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07864_ _02865_ register_file\[6\]\[24\] _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09603_ _04912_ _04914_ _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07795_ register_file\[3\]\[23\] _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09534_ _04576_ register_file\[7\]\[14\] _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13462__A1 _07572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__A2 register_file\[18\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09465_ _04712_ register_file\[12\]\[13\] _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08416_ _03741_ _03743_ _03436_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13214__A1 _07619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09396_ _04710_ register_file\[17\]\[12\] _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09969__A1 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08347_ _01176_ _03673_ _03675_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08278_ _03588_ _03607_ _03303_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11528__A1 _06558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15684__CLK clknet_leaf_70_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10240_ _05275_ register_file\[15\]\[24\] _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10235__B _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10200__A1 _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_254_clk clknet_5_16__leaf_clk clknet_leaf_254_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_161_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10171_ _05273_ register_file\[26\]\[23\] _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08944__A2 register_file\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10751__A2 register_file\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15317__I _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13930_ register_file\[5\]\[3\] _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11700__A1 _06663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10503__A2 register_file\[25\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13861_ _01377_ _01378_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15600_ _03077_ _03097_ _02762_ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15442__A2 register_file\[13\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12812_ _07241_ _07360_ _07367_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16580_ _00968_ clknet_leaf_57_clk register_file\[9\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12256__A2 register_file\[31\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13453__A1 _07562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13792_ _01310_ _01063_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15531_ _02857_ register_file\[14\]\[22\] _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12743_ _07313_ _07326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15462_ _02954_ _02961_ _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12674_ _07231_ _07279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13205__A1 _07612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12008__A2 _06854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08880__A1 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10019__A1 _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14413_ _01755_ register_file\[22\]\[9\] _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14891__I _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11625_ _06613_ register_file\[10\]\[15\] _06617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13756__A2 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15393_ _02892_ _02808_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11767__A1 _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14344_ _01682_ register_file\[11\]\[8\] _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11556_ _06553_ _06575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_102_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10507_ _05609_ register_file\[27\]\[28\] _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14275_ register_file\[4\]\[7\] _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_155_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11487_ _06429_ _06527_ _06533_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16014_ _00402_ clknet_leaf_246_clk register_file\[6\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09188__A2 register_file\[13\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13226_ _07576_ _07622_ _07627_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14181__A2 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10438_ _05672_ register_file\[13\]\[27\] _05738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12192__A1 _06969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_245_clk clknet_5_17__leaf_clk clknet_leaf_245_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13157_ _07502_ _07584_ _07587_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _05667_ _05669_ _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12108_ _06649_ _06912_ _06919_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13088_ _06084_ _07538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12039_ _06865_ _06878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08699__A1 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13692__A1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15433__A2 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12247__A2 _07000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09112__A2 register_file\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15729_ _00117_ clknet_leaf_166_clk register_file\[27\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13995__A2 _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09250_ _04565_ _04566_ _04567_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08201_ _03459_ register_file\[1\]\[28\] _01198_ _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09181_ _04499_ register_file\[3\]\[8\] _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11758__A1 _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08132_ _03443_ _03463_ _03303_ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08623__A1 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10430__A1 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08063_ _03063_ register_file\[19\]\[27\] _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09179__A2 register_file\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14172__A2 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_242_clk_I clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11930__A1 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08965_ _04283_ _04286_ _03914_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11665__I _06639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14041__I _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07916_ _03084_ register_file\[18\]\[25\] _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12486__A2 register_file\[23\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_257_clk_I clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08896_ _03875_ _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__13683__A1 _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input24_I new_value[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10497__A1 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07847_ _03181_ register_file\[8\]\[24\] _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07778_ _02857_ register_file\[14\]\[23\] _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13435__A1 _07749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10249__A1 _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09517_ _04830_ register_file\[10\]\[13\] _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16482__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11997__A1 _06698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09448_ _04753_ _04762_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08862__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09379_ _04685_ _04694_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08923__B _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11749__A1 _06698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11410_ _06431_ _06486_ _06487_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12390_ _06980_ _07098_ _07101_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08614__A1 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12410__A2 _07112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10421__A1 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10744__I _06036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11341_ _06368_ register_file\[19\]\[31\] _06445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08090__A2 _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output92_I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10972__A2 _06206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14060_ _01575_ _01488_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11272_ _06391_ register_file\[19\]\[10\] _06397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12174__A1 _06716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13011_ _07281_ _07480_ _07486_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10223_ _05525_ register_file\[22\]\[24\] _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13910__A2 _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11921__A1 _06803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _05254_ register_file\[16\]\[23\] _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14962_ _02466_ _02467_ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12477__A2 register_file\[23\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10085_ _05190_ register_file\[26\]\[22\] _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09342__A2 register_file\[21\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10488__A1 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13913_ _01125_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14893_ _01559_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13844_ _01357_ _01362_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12229__A2 register_file\[31\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13426__A1 _07536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10919__I _06169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16563_ _00951_ clknet_leaf_179_clk register_file\[29\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13775_ _01015_ register_file\[19\]\[2\] _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10987_ _06217_ _06218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15179__A1 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15514_ _03006_ _03012_ _02924_ _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12726_ _07314_ register_file\[20\]\[1\] _07316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16494_ _00882_ clknet_leaf_188_clk register_file\[15\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15445_ _01693_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12657_ _07234_ _07267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15510__I _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11608_ _06606_ register_file\[10\]\[8\] _06607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15376_ _01175_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12401__A2 register_file\[24\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12588_ _07219_ register_file\[22\]\[23\] _07220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16205__CLK clknet_leaf_138_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14327_ _01083_ _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11539_ _06545_ _06565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08081__A2 register_file\[26\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14154__A2 _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14258_ _01768_ _01771_ _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12165__A1 _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_218_clk clknet_5_23__leaf_clk clknet_leaf_218_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13209_ _07612_ register_file\[15\]\[22\] _07618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08908__A2 register_file\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14189_ register_file\[4\]\[6\] _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11912__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16355__CLK clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08750_ _03908_ register_file\[31\]\[2\] _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12468__A2 _07146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09333__A2 register_file\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08681_ _04004_ _04005_ _04006_ _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13914__B _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13417__A1 _07526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10829__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09097__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13968__A2 register_file\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14090__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09302_ _04348_ register_file\[27\]\[10\] _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11979__A1 _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08844__A1 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09233_ _04348_ register_file\[19\]\[9\] _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09164_ _04346_ register_file\[26\]\[8\] _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14393__A2 register_file\[30\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15590__A1 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08115_ _03444_ _03446_ _03369_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10403__A1 _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08072__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09095_ _03770_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_181_clk_I clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10954__A2 register_file\[2\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08034__I register_file\[7\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08046_ _03378_ _03210_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12156__A1 _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_209_clk clknet_5_23__leaf_clk clknet_leaf_209_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_150_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_61_clk_I clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14696__A3 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08969__I _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09021__A1 _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09997_ _05303_ register_file\[2\]\[20\] _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_196_clk_I clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08948_ _04054_ register_file\[31\]\[5\] _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12459__A2 register_file\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_76_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _04197_ _04200_ _04201_ _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11131__A2 register_file\[27\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10910_ _06170_ register_file\[2\]\[1\] _06172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11890_ _06672_ _06785_ _06788_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10739__I _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10841_ _06115_ _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13959__A2 register_file\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09088__A1 _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14081__A1 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13560_ _01080_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ _06059_ _06060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_158_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12631__A2 register_file\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_134_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12511_ _07021_ _07167_ _07173_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10642__A1 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09749__B _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13491_ _01007_ _01011_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15230_ _02651_ register_file\[20\]\[19\] _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_clk_I clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12442_ _07032_ _07126_ _07131_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14384__A2 register_file\[27\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15581__A1 _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12395__A1 _06985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11198__A2 _06344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15161_ _02663_ _02331_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09260__A1 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12373_ _06958_ _07088_ _07091_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08063__A2 register_file\[19\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10945__A2 register_file\[2\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14112_ _01369_ register_file\[1\]\[5\] _01371_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14136__A2 register_file\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16378__CLK clknet_leaf_255_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11324_ _06431_ _06432_ _06433_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15092_ _02589_ _02595_ _02508_ _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_158_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07810__A2 register_file\[19\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12147__A1 _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_29_clk_I clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14043_ _01074_ _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__A1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11255_ _06378_ register_file\[19\]\[5\] _06385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10206_ _05306_ register_file\[1\]\[23\] _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11186_ _06082_ _06337_ _06340_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10137_ _05306_ register_file\[1\]\[22\] _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15994_ _00382_ clknet_leaf_252_clk register_file\[7\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10068_ _05173_ register_file\[3\]\[21\] _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14945_ _02450_ register_file\[6\]\[15\] _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11122__A2 register_file\[27\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08828__B _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14876_ _02045_ _02380_ _02382_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07877__A2 register_file\[2\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12870__A2 _07398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10881__A1 _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13827_ _01342_ _01343_ _01345_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14611__A3 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16546_ _00934_ clknet_leaf_19_clk register_file\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08826__A1 _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13758_ _01277_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_62_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12709_ _07302_ _07296_ _07303_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12864__I _07369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16477_ _00865_ clknet_leaf_301_clk register_file\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13689_ _01019_ register_file\[18\]\[1\] _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15572__A1 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15428_ _02764_ register_file\[8\]\[21\] _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11189__A2 _06337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12386__A1 _06974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15359_ _02859_ register_file\[15\]\[20\] _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09251__A1 _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10936__A2 _06185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12138__A1 _06679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09920_ _03879_ _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09394__B _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15745__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12689__A2 _07284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09851_ _05158_ _05159_ _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09554__A2 register_file\[13\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08357__A3 _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08802_ _04125_ register_file\[24\]\[3\] _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09782_ _05089_ _05091_ _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08733_ _04051_ _04056_ _04057_ _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11113__A2 _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12310__A1 _06980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08664_ _03987_ _03989_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12861__A2 _07391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10872__A1 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14063__A1 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08595_ _03776_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09490__A1 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08293__A2 register_file\[23\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07868__I _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09216_ _04257_ register_file\[22\]\[9\] _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16520__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12377__A1 _06967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09147_ _04259_ register_file\[23\]\[8\] _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09078_ _04259_ register_file\[23\]\[7\] _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12129__A1 _06926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ _03276_ register_file\[15\]\[26\] _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11040_ _06247_ register_file\[28\]\[20\] _06251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11352__A2 register_file\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output55_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15094__A3 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12991_ _07470_ register_file\[17\]\[11\] _07475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15325__I _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12301__A1 _07046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14730_ _02236_ _01901_ _02237_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14841__A3 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11942_ _06818_ register_file\[5\]\[1\] _06820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07859__A2 register_file\[14\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14661_ _02169_ register_file\[20\]\[12\] _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11873_ _06774_ register_file\[6\]\[5\] _06779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16050__CLK clknet_leaf_230_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16400_ _00788_ clknet_leaf_160_clk register_file\[18\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13612_ _01132_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10824_ net19 _06102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14592_ _02101_ register_file\[11\]\[11\] _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15618__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12604__A2 _07186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13801__A1 _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16331_ _00719_ clknet_leaf_137_clk register_file\[20\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12684__I _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13543_ _01061_ _01063_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10755_ _06045_ _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09481__A1 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08284__A2 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16262_ _00650_ clknet_leaf_91_clk register_file\[22\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10091__A2 register_file\[29\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13474_ _00994_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14357__A2 register_file\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15554__A1 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10686_ _03901_ register_file\[16\]\[31\] _05982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15213_ _02714_ _02715_ _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12425_ _07116_ register_file\[24\]\[22\] _07122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16193_ _00581_ clknet_leaf_70_clk register_file\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09233__A1 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10918__A2 _06168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11040__A1 _06247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15144_ _02646_ register_file\[19\]\[18\] _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09784__A2 register_file\[31\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12356_ _07026_ _07078_ _07080_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11307_ _06419_ _06420_ _06421_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11591__A2 _06592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10932__I _06177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15075_ _02578_ _02331_ _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12287_ _06317_ _03794_ _07038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_45_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14026_ _01177_ _01540_ _01542_ _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11238_ _06366_ _06369_ _06372_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11343__A2 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12540__A1 _06969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_27__f_clk clknet_3_6_0_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_150_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11169_ _06326_ register_file\[13\]\[5\] _06331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12859__I _07358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15977_ _00365_ clknet_leaf_291_clk register_file\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11763__I _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14928_ _02433_ _02272_ _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12843__A2 register_file\[1\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10854__A1 _06109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14859_ _02358_ _02365_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08380_ register_file\[11\]\[31\] _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16543__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10606__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16529_ _00917_ clknet_leaf_172_clk register_file\[14\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09472__A1 _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10082__A2 register_file\[25\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09001_ _04318_ _04321_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12359__A1 _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08027__A2 register_file\[14\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11003__I _06228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13020__A2 register_file\[17\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10909__A2 _06168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11031__A1 _06100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09775__A2 register_file\[7\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11938__I _06814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11582__A2 _06546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10842__I _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13859__A1 _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09903_ _05203_ _05210_ _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09527__A2 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09834_ _05139_ _05142_ _04002_ _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09852__B _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09765_ _05073_ _05074_ _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16073__CLK clknet_leaf_289_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13087__A2 _07532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11098__A1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ _04039_ _04040_ _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09696_ _04937_ register_file\[30\]\[16\] _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12834__A2 _07377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10845__A1 _06117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08647_ _03969_ _03972_ _03856_ _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14587__A2 register_file\[9\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08578_ _03904_ _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12598__A1 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_165_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08266__A2 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15910__CLK clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15536__A1 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10540_ _05825_ _05838_ _05839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_195_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10471_ _05769_ _05770_ _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13011__A2 _07480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08931__B _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12210_ _06982_ _06976_ _06984_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13190_ _07605_ register_file\[15\]\[14\] _07607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12770__A1 _07340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11573__A2 register_file\[11\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12141_ _06933_ register_file\[3\]\[17\] _06939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14511__A2 register_file\[12\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12072_ _02955_ _06895_ _06897_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12522__A1 _07032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11023_ _06240_ register_file\[28\]\[13\] _06241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15900_ _00288_ clknet_leaf_283_clk register_file\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16416__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15831_ _00219_ clknet_leaf_219_clk register_file\[26\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11089__A1 _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15762_ _00150_ clknet_leaf_177_clk register_file\[13\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12974_ _07244_ _07456_ _07464_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12825__A2 _07370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16566__CLK clknet_leaf_215_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14713_ _02212_ _02221_ _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10199__I _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11925_ _06803_ register_file\[6\]\[27\] _06809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14027__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15693_ _00081_ clknet_leaf_148_clk register_file\[28\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14578__A2 register_file\[22\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14644_ _01904_ register_file\[30\]\[12\] _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11856_ _06766_ _06767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12589__A1 _07018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10807_ _06086_ _06074_ _06088_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10927__I _06169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14575_ _01751_ register_file\[20\]\[11\] _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11787_ _06726_ register_file\[7\]\[3\] _06727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13250__A2 _07642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11261__A1 _06378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16314_ _00702_ clknet_leaf_270_clk register_file\[21\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13526_ _01037_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10738_ _06031_ _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16245_ _00633_ clknet_leaf_183_clk register_file\[23\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09206__A1 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13457_ _07763_ register_file\[9\]\[25\] _07767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13002__A2 _07480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10669_ _05961_ _05964_ _04037_ _05965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12408_ _07097_ _07112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11013__A1 _06233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16176_ _00564_ clknet_leaf_154_clk register_file\[25\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13388_ _07578_ _07682_ _07724_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput106 net106 rS[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_114_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12761__A1 _07333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11564__A2 register_file\[11\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12339_ _07009_ _07064_ _07070_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15127_ register_file\[3\]\[17\] _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09509__A2 register_file\[31\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15058_ _02561_ _02228_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11316__A2 register_file\[19\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13973__I _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12513__A1 _07171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16096__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14009_ _01152_ register_file\[6\]\[4\] _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_29_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07880_ _02877_ _03212_ _03214_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07971__I _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13069__A2 register_file\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14266__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09550_ _04661_ register_file\[30\]\[14\] _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08501_ _03827_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10827__A1 _06087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09481_ _04729_ register_file\[16\]\[13\] _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14018__A1 _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15933__CLK clknet_leaf_307_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08432_ _03740_ _03759_ _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14569__A2 _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10837__I _06112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08363_ _03685_ _03690_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09445__A1 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13241__A2 _07632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15518__A1 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08294_ _03621_ _01094_ _03622_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10058__B _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11004__A1 _06225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11668__I _06642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12752__A1 _07262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11555__A2 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16439__CLK clknet_leaf_204_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14044__I _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12504__A1 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11307__A2 _06420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08184__A1 _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16589__CLK clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_10__f_clk clknet_3_2_0_clk clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09817_ _04855_ register_file\[7\]\[18\] _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09748_ _05056_ _05057_ _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12807__A2 _07360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10818__A1 _06095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09679_ _04988_ _04989_ _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14009__A1 _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11710_ _06663_ register_file\[8\]\[12\] _06673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11491__A1 _06531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10294__A2 _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12690_ _06129_ _07290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09601__I _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11641_ _06620_ register_file\[10\]\[22\] _06626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09436__A1 _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10747__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13123__I _07503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10046__A2 register_file\[14\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15509__A1 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14360_ _01870_ _01872_ _01702_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11243__A1 _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11572_ _06434_ _06582_ _06584_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13311_ _06316_ _03815_ _07678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07998__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12991__A1 _07470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10523_ _05695_ register_file\[31\]\[28\] _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11794__A2 _06730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput19 new_value[17] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14291_ _01795_ _01804_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12962__I _07454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16030_ _00418_ clknet_leaf_298_clk register_file\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13242_ _07633_ _07638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09739__A2 register_file\[10\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10454_ _05751_ _05753_ _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14732__A2 register_file\[31\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11546__A2 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13173_ _07590_ register_file\[15\]\[7\] _07597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10385_ _05416_ register_file\[14\]\[26\] _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12124_ _06921_ _06929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14496__A1 _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13299__A2 register_file\[14\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12055_ _02372_ _06881_ _06887_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08175__A1 _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11006_ _06225_ register_file\[28\]\[6\] _06231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07922__A1 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15956__CLK clknet_leaf_221_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15814_ _00202_ clknet_leaf_107_clk register_file\[26\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15745_ _00133_ clknet_leaf_53_clk register_file\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09675__A1 _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12957_ _07407_ register_file\[18\]\[31\] _07453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11482__A1 _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11908_ _06777_ _06799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15676_ _00064_ clknet_leaf_36_clk register_file\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12888_ _07410_ register_file\[18\]\[2\] _07413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14627_ _02135_ _02136_ _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11839_ _06701_ _06751_ _06757_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10037__A2 register_file\[30\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09978__A2 register_file\[7\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08127__I _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14558_ _01986_ register_file\[29\]\[11\] _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14971__A2 register_file\[25\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14573__B _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12982__A1 _07252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11785__A2 _06720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13509_ _01029_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14489_ _01746_ register_file\[19\]\[10\] _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16228_ _00616_ clknet_leaf_77_clk register_file\[23\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14723__A2 register_file\[27\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11488__I _06505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12734__A1 _07244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16159_ _00547_ clknet_leaf_17_clk register_file\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_192_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08981_ _04233_ register_file\[7\]\[6\] _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07932_ _03265_ _03104_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07863_ _03190_ _03197_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14239__A1 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09602_ _04913_ register_file\[27\]\[15\] _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12112__I _06921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07794_ _02964_ register_file\[2\]\[23\] _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_3_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09533_ _04781_ register_file\[6\]\[14\] _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11951__I _06817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13462__A2 _07766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11473__A1 _06414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09464_ _04710_ register_file\[13\]\[13\] _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16111__CLK clknet_leaf_190_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08415_ _03742_ _01097_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09395_ _03766_ _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09418__A1 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14411__A1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13214__A2 register_file\[15\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08346_ _03674_ _01156_ _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11225__A1 _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09969__A2 register_file\[27\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12973__A1 _07462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16261__CLK clknet_leaf_75_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09577__B _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08277_ _03599_ _03606_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12725__A1 _07230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10200__A2 register_file\[23\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _05472_ _05473_ _05474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14478__A1 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08157__A1 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13150__A1 _07580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10251__B _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07904__A1 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11700__A2 register_file\[8\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13860_ _01000_ register_file\[17\]\[3\] _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14658__B _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12811_ _07366_ register_file\[1\]\[3\] _07367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09657__A1 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13791_ _01306_ _01309_ _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08656__B _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13453__A2 _07759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15530_ _03025_ _03026_ _03028_ _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12742_ _07252_ _07322_ _07325_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12673_ _06107_ _07278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15461_ _02956_ _02959_ _02960_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13205__A2 register_file\[15\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_190_clk clknet_5_25__leaf_clk clknet_leaf_190_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08880__A2 register_file\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14412_ _01922_ _01840_ _01923_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10019__A2 register_file\[19\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11624_ _06601_ _06616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15392_ _02890_ _02891_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13788__I _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11767__A2 register_file\[8\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12964__A1 _07458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11555_ _06417_ _06568_ _06574_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14343_ _01854_ _01855_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10506_ _05607_ register_file\[26\]\[28\] _05805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14274_ _01784_ _01787_ _01702_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11486_ _06531_ register_file\[12\]\[24\] _06533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16013_ _00401_ clknet_leaf_247_clk register_file\[6\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13225_ _07583_ register_file\[15\]\[29\] _07627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10437_ _05733_ _05736_ _05268_ _05737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12192__A2 _06961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13156_ _07586_ register_file\[15\]\[0\] _07587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10368_ _05668_ register_file\[7\]\[26\] _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15508__I _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12107_ _06918_ register_file\[3\]\[3\] _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13087_ _07536_ _07532_ _07537_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10299_ _05334_ register_file\[11\]\[25\] _05601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13141__A1 _07574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12038_ _01789_ _06874_ _06877_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09896__A1 _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08699__A2 register_file\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09648__A1 _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14641__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13989_ _01505_ _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15728_ _00116_ clknet_leaf_166_clk register_file\[27\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11455__A1 _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08320__A1 _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15659_ _00047_ clknet_leaf_141_clk register_file\[2\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16284__CLK clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_181_clk clknet_5_28__leaf_clk clknet_leaf_181_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08871__A2 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08200_ _03294_ _03528_ _03530_ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_178_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11207__A1 _06348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09180_ _03919_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13747__A3 _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11758__A2 register_file\[8\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08131_ _03454_ _03462_ _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12955__A1 _07407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09820__A1 _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08062_ _03393_ _02978_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10430__A2 register_file\[9\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13380__A1 _07570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10194__A1 _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11946__I _06817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11930__A2 _06806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14322__I _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08964_ _04284_ _04285_ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08139__A1 _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13132__A1 _07567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07915_ _02998_ register_file\[19\]\[25\] _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08895_ _04216_ _04217_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14880__A1 _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13683__A2 register_file\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07846_ _01079_ _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10497__A2 register_file\[4\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11694__A1 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input17_I new_value[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07777_ _03111_ _03026_ _03112_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_77_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14632__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11681__I _06045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09516_ _04145_ _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11446__A1 _06388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10249__A2 register_file\[7\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13986__A3 _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09447_ _04758_ _04761_ _04486_ _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11997__A2 _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_172_clk clknet_5_29__leaf_clk clknet_leaf_172_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09378_ _04688_ _04693_ _03894_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14935__A2 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15651__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11749__A2 _06692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12946__A1 _07295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08329_ _03657_ register_file\[15\]\[30\] _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15102__B _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11340_ _06163_ _06444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_192_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16007__CLK clknet_leaf_297_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11271_ _06383_ _06396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12017__I _06863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15360__A2 _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13010_ _07484_ register_file\[17\]\[19\] _07486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output85_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10222_ _03867_ _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12174__A2 _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_8__f_clk clknet_3_2_0_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11856__I _06766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14232__I _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _05252_ register_file\[17\]\[23\] _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10760__I _06049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16157__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10084_ _05387_ _05388_ _05389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14961_ _02217_ register_file\[1\]\[15\] _02218_ _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13912_ _01249_ register_file\[10\]\[3\] _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14892_ _02397_ register_file\[26\]\[15\] _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12687__I _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13843_ _01359_ _01361_ _01273_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13426__A2 _07745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11437__A1 _06502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16562_ _00950_ clknet_leaf_180_clk register_file\[29\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10986_ _04077_ _06216_ _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13774_ _01291_ _01292_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08302__A1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15513_ _03008_ _03009_ _03011_ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_188_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12725_ _07230_ _07312_ _07315_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16493_ _00881_ clknet_leaf_125_clk register_file\[15\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15179__A2 register_file\[8\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08853__A2 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09996__I _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_302_clk_I clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15444_ _02857_ register_file\[14\]\[21\] _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12656_ _06085_ _07266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10660__A2 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12937__A1 _07436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11607_ _06593_ _06606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14407__I _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12587_ _07182_ _07219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15375_ _02875_ _02793_ _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14326_ _01751_ register_file\[20\]\[8\] _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11538_ _06400_ _06561_ _06564_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11469_ _06517_ register_file\[12\]\[17\] _06523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14257_ _01769_ _01770_ _01431_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13362__A1 _07708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13208_ _07558_ _07615_ _07617_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10176__A1 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14188_ _01699_ _01701_ _01702_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13901__A3 _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11766__I _06155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11912__A2 _06799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13139_ _06150_ _07574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13114__A1 _07551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I addrS[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09680__B _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11676__A1 _06647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08680_ _03923_ register_file\[1\]\[1\] _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15406__A3 _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13417__A2 _07738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11428__A1 _06498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09097__A2 register_file\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15674__CLK clknet_leaf_257_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09301_ _04346_ register_file\[26\]\[10\] _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14090__A2 register_file\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_154_clk clknet_5_30__leaf_clk clknet_leaf_154_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10100__A1 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08844__A2 register_file\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09232_ _04346_ register_file\[18\]\[9\] _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14917__A2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12928__A1 _07436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09163_ _04480_ _04481_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15590__A2 register_file\[20\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_10__f_clk_I clknet_3_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08114_ _03445_ _01167_ _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09094_ _04413_ register_file\[5\]\[7\] _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10066__B _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ _03370_ _03377_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13353__A1 _07701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12156__A2 register_file\[3\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15148__I _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09996_ _03779_ _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08947_ _04052_ register_file\[30\]\[5\] _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14853__A1 _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08878_ _03894_ _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07829_ _03162_ _03163_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10840_ net23 _06115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11419__A1 _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10771_ _06058_ _06059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_145_clk clknet_5_27__leaf_clk clknet_leaf_145_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12510_ _07171_ register_file\[23\]\[24\] _07173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13490_ _01010_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12919__A1 _07269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12441_ _07087_ register_file\[24\]\[29\] _07131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14227__I _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10755__I _06045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15581__A2 register_file\[17\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12395__A2 _07098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15160_ _02661_ _02662_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12372_ _07090_ register_file\[24\]\[0\] _07091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09260__A2 register_file\[31\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14111_ _01623_ _01624_ _01626_ _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11323_ _06427_ register_file\[19\]\[25\] _06433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15091_ _02591_ _02592_ _02594_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12970__I _07457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13344__A1 _07534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12147__A2 _06936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11254_ _06383_ _06384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_14042_ _01557_ register_file\[26\]\[5\] _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11586__I _06590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13895__A2 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10205_ _05508_ register_file\[3\]\[23\] _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11185_ _06334_ register_file\[13\]\[12\] _06340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10136_ _05173_ register_file\[3\]\[22\] _05441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14897__I _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15993_ _00381_ clknet_leaf_243_clk register_file\[7\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14844__A1 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13647__A2 _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10067_ _05303_ register_file\[2\]\[21\] _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14944_ _01178_ _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11658__A1 _06440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15697__CLK clknet_leaf_166_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14875_ _02381_ _02300_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13826_ _01344_ register_file\[13\]\[2\] _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10881__A2 register_file\[30\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_241_clk_I clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16545_ _00933_ clknet_leaf_18_clk register_file\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_136_clk clknet_5_26__leaf_clk clknet_leaf_136_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13757_ _01178_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10969_ _06203_ register_file\[2\]\[25\] _06207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12708_ _07232_ register_file\[21\]\[28\] _07303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11830__A1 _06691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16476_ _00864_ clknet_leaf_282_clk register_file\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15021__A1 _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13688_ _01015_ register_file\[19\]\[1\] _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15427_ _02907_ _02926_ _02762_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12639_ _06063_ _07254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15572__A2 register_file\[29\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13041__I _07503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12386__A2 _07098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_256_clk_I clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16322__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15358_ _01455_ _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09251__A2 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14309_ _01478_ register_file\[30\]\[8\] _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12880__I _07406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15289_ _02788_ _02790_ _02544_ _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_171_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12138__A2 _06936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10149__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16472__CLK clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ _05025_ register_file\[19\]\[18\] _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11897__A1 _06789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08762__A1 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08801_ _04124_ _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09781_ _05090_ register_file\[28\]\[17\] _05091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14835__A1 _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08732_ _03913_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11649__A1 _06627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12310__A2 _07050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08663_ _03988_ register_file\[23\]\[1\] _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10321__A1 _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13216__I _07593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10872__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08594_ _03920_ register_file\[3\]\[0\] _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14063__A2 register_file\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_209_clk_I clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_127_clk clknet_5_25__leaf_clk clknet_leaf_127_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_41_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13810__A2 _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08754__B _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11821__A1 _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09490__A2 register_file\[22\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09215_ _04531_ _04532_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15563__A2 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09146_ _04257_ register_file\[22\]\[8\] _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12377__A2 _07088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14491__B _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09077_ _04257_ register_file\[22\]\[7\] _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12129__A2 register_file\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13326__A1 _07516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08028_ _01693_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11888__A1 _06670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15079__A1 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09979_ _05284_ _05285_ _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10560__A1 _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15606__I _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12990_ _07259_ _07473_ _07474_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output48_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11941_ _06638_ _06816_ _06819_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10312__A1 _05596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14660_ _01318_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11872_ _06777_ _06778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13611_ _01034_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10823_ _06100_ _06096_ _06101_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14591_ _01681_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16330_ _00718_ clknet_leaf_99_clk register_file\[20\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11812__A1 _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13542_ _01062_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16345__CLK clknet_leaf_196_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10754_ _06044_ _06045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16261_ _00649_ clknet_leaf_75_clk register_file\[22\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13473_ _00993_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15554__A2 register_file\[1\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10685_ _03898_ register_file\[17\]\[31\] _05981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15212_ _01155_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12424_ _07014_ _07119_ _07121_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16192_ _00580_ clknet_leaf_11_clk register_file\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09233__A2 register_file\[19\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15143_ _01068_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16495__CLK clknet_leaf_188_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11040__A2 register_file\[28\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12355_ _07075_ register_file\[25\]\[26\] _07080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08992__A1 _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13317__A1 _07502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11306_ _06415_ register_file\[19\]\[20\] _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15074_ _02575_ _02577_ _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12286_ _07036_ _06963_ _07037_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14025_ _01541_ _01456_ _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11237_ _06371_ register_file\[19\]\[0\] _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12540__A2 _07184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11168_ _06329_ _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14817__A1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10119_ _05423_ register_file\[13\]\[22\] _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14420__I _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11099_ _06073_ _06286_ _06287_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15976_ _00364_ clknet_leaf_297_clk register_file\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14927_ _02432_ _02270_ _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10303__A1 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_180_clk_I clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14858_ _02361_ _02364_ _02030_ _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10854__A2 register_file\[30\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15242__A1 _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13809_ _01327_ register_file\[31\]\[2\] _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_109_clk clknet_5_12__leaf_clk clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_60_clk_I clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14789_ _02296_ _01961_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07969__I _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16528_ _00916_ clknet_leaf_173_clk register_file\[14\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11803__A1 _06665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09472__A2 register_file\[25\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10609__B _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_195_clk_I clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16459_ _00847_ clknet_leaf_130_clk register_file\[16\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15712__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09000_ _04320_ register_file\[19\]\[6\] _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12359__A2 register_file\[25\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_7_0_clk clknet_0_clk clknet_3_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_75_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11031__A2 _06243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13308__A1 _07578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08983__A1 _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10790__A1 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13859__A2 register_file\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09902_ _05206_ _05209_ _04553_ _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14520__A3 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08735__A1 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09833_ _05140_ _05141_ _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10542__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09764_ _04939_ register_file\[23\]\[17\] _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_13_clk_I clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15481__A1 _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14284__A2 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08715_ _03967_ register_file\[12\]\[2\] _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11098__A2 register_file\[27\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12295__A1 _06965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09695_ _05003_ _05005_ _05006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_148_clk_I clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10845__A2 _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08646_ _03970_ _03971_ _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12047__A1 _06878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_28_clk_I clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08577_ _03806_ _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_161_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12598__A2 _07222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13795__A1 _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15536__A2 register_file\[6\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10470_ _05503_ register_file\[27\]\[27\] _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09129_ _04446_ _04447_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07777__A2 _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12140_ _06682_ _06936_ _06938_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08974__A1 _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12770__A2 register_file\[20\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08503__I _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12071_ _06892_ net24 _06897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11022_ _06220_ _06240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12522__A2 _07174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15830_ _00218_ clknet_leaf_219_clk register_file\[26\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15472__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15761_ _00149_ clknet_leaf_173_clk register_file\[13\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11089__A2 _06279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12286__A1 _07036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12973_ _07462_ register_file\[17\]\[4\] _07464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14712_ _02220_ _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11924_ _06706_ _06806_ _06808_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15692_ _00080_ clknet_leaf_134_clk register_file\[28\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14643_ _02150_ _01901_ _02151_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11855_ _06024_ _03913_ _06766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12589__A2 _07215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10806_ _06087_ register_file\[30\]\[13\] _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14574_ _02080_ _02083_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11786_ _06721_ _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08257__A3 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16313_ _00701_ clknet_leaf_194_clk register_file\[21\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13525_ _01045_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11261__A2 register_file\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10737_ net22 _06031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11104__I _06270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16244_ _00632_ clknet_leaf_181_clk register_file\[23\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13456_ _07737_ _07766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_103_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10668_ _05962_ _05963_ _05964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12407_ _06997_ _07105_ _07111_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16175_ _00563_ clknet_leaf_144_clk register_file\[25\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12210__A1 _06982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11013__A2 register_file\[28\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13387_ _07679_ register_file\[29\]\[30\] _07724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10599_ _05896_ _05643_ _05897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput107 net107 rS[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__12761__A2 register_file\[20\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15126_ _02548_ register_file\[2\]\[17\] _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12338_ _07068_ register_file\[25\]\[19\] _07070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15057_ _02560_ _02393_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09953__B _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12269_ _06143_ _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08717__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12513__A2 register_file\[23\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14008_ _01517_ _01524_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08193__A2 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16510__CLK clknet_leaf_305_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12277__A1 _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15959_ _00347_ clknet_leaf_239_clk register_file\[8\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08500_ _03778_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10827__A2 register_file\[30\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09480_ _04727_ register_file\[17\]\[13\] _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15215__A1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14018__A2 _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12029__A1 _06870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08431_ _03749_ _03758_ _01011_ _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_145_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08362_ _03687_ _03689_ _01035_ _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09445__A2 register_file\[27\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08293_ _03320_ register_file\[23\]\[30\] _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15518__A2 register_file\[9\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10853__I _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11004__A2 register_file\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12752__A2 _07329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10074__B _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10763__A1 _06042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08420__A3 _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16040__CLK clknet_leaf_296_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12504__A2 _07167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13701__A1 _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10515__A1 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11684__I _06049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09381__A1 _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09816_ _04853_ register_file\[6\]\[18\] _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09154__I _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16190__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07931__A2 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09747_ _04855_ register_file\[27\]\[17\] _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12268__A1 _07023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15758__CLK clknet_leaf_148_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10818__A2 _06096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09678_ _04855_ register_file\[23\]\[16\] _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14009__A2 register_file\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08629_ _03953_ _03954_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13768__A1 _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11640_ _06422_ _06623_ _06625_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08239__A3 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15509__A2 register_file\[30\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12440__A1 _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11571_ _06579_ register_file\[11\]\[26\] _06584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13310_ _07580_ _07634_ _07677_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07998__A2 register_file\[26\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12991__A2 register_file\[17\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10522_ _05693_ register_file\[30\]\[28\] _05821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14290_ _01803_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11859__I _06769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14193__A1 _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10453_ _05752_ register_file\[7\]\[27\] _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13241_ _07511_ _07632_ _07637_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__A1 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13940__A1 _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13172_ _07522_ _07594_ _07596_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10384_ _05683_ _05684_ _05685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08411__A3 _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12123_ _06665_ _06922_ _06928_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14496__A2 register_file\[22\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12054_ _06885_ net16 _06887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10506__A1 _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11594__I _06593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11005_ _06050_ _06229_ _06230_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14248__A2 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15813_ _00201_ clknet_leaf_64_clk register_file\[26\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14799__A3 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09124__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09999__I _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15744_ _00132_ clknet_leaf_4_clk register_file\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12956_ _07306_ _07410_ _07452_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09675__A2 register_file\[20\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11907_ _06689_ _06792_ _06798_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11482__A2 _06527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15675_ _00063_ clknet_leaf_284_clk register_file\[2\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12887_ _07237_ _07408_ _07412_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13314__I _07678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13759__A1 _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14626_ _01800_ register_file\[1\]\[11\] _01801_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11838_ _06755_ register_file\[7\]\[24\] _06757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10159__B _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12431__A1 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14557_ _01818_ register_file\[28\]\[11\] _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11769_ _06159_ _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_clk clknet_5_13__leaf_clk clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08852__B _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13508_ _00992_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07989__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12982__A2 _07466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14488_ _01998_ _01832_ _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10993__A1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11769__I _06159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16227_ _00615_ clknet_leaf_78_clk register_file\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14184__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13439_ _07726_ _07756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08938__A1 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12734__A2 _07312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16158_ _00546_ clknet_leaf_24_clk register_file\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10745__A1 _06029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08402__A3 _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15109_ _02442_ register_file\[14\]\[17\] _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16089_ _00477_ clknet_leaf_248_clk register_file\[4\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08980_ _04090_ register_file\[6\]\[6\] _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14487__A2 _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07931_ _03264_ _03102_ _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12498__A1 _07164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09363__A1 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15900__CLK clknet_leaf_283_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07862_ _03193_ _03196_ _02862_ _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11170__A1 _06050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14239__A2 register_file\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09601_ _03785_ _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07913__A2 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07793_ _03128_ _02793_ _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09115__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09532_ _02374_ _03763_ _04844_ _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13998__A1 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10848__I _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09463_ _04744_ _04777_ _04641_ net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11473__A2 _06520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08414_ register_file\[17\]\[31\] _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09394_ _04678_ _04709_ _04641_ net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09418__A2 register_file\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14411__A2 register_file\[21\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12422__A1 _07011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08345_ register_file\[3\]\[30\] _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__16406__CLK clknet_leaf_214_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08762__B _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ _03605_ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12973__A2 register_file\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14175__A1 _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14714__A3 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08929__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12725__A2 _07312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10736__A1 _06021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14478__A2 register_file\[30\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12489__A1 _07157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98_clk clknet_5_15__leaf_clk clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09354__A1 _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13150__A2 _07507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12303__I _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11161__A1 _06037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07904__A2 register_file\[30\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12810_ _07361_ _07366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13790_ _01308_ register_file\[25\]\[2\] _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12741_ _07318_ register_file\[20\]\[7\] _07325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10758__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12661__A1 _07267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15460_ _01034_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12672_ _07276_ _07272_ _07277_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14411_ _01841_ register_file\[21\]\[9\] _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11623_ _06405_ _06609_ _06615_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16086__CLK clknet_leaf_234_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12413__A1 _07109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15391_ _02805_ register_file\[17\]\[21\] _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_22_clk clknet_5_2__leaf_clk clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14953__A3 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14342_ _01426_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11554_ _06572_ register_file\[11\]\[19\] _06574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10707__B _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10975__A1 _06167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10505_ _05802_ _05803_ _05804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07840__A1 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14273_ _01785_ _01786_ _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11485_ _06426_ _06527_ _06532_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16012_ _00400_ clknet_leaf_249_clk register_file\[6\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13224_ _07574_ _07622_ _07626_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10436_ _05734_ _05735_ _05736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10727__A1 _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08396__A2 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13155_ _07585_ _07586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15923__CLK clknet_leaf_213_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10367_ _04319_ _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12106_ _06913_ _06918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13086_ _07527_ register_file\[16\]\[12\] _07537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10298_ _05332_ register_file\[10\]\[25\] _05600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_89_clk clknet_5_14__leaf_clk clknet_leaf_89_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08148__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13141__A2 _07568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12037_ _06870_ net40 _06877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15418__A1 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09896__A2 register_file\[17\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13988_ net10 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09648__A2 register_file\[21\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14641__A2 register_file\[28\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15727_ _00115_ clknet_5_27__leaf_clk register_file\[27\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12652__A1 _07262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12939_ _07406_ _07443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11455__A2 register_file\[12\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16429__CLK clknet_leaf_142_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13044__I _07506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15658_ _00046_ clknet_leaf_94_clk register_file\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15197__A3 _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14609_ _02118_ _01786_ _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12404__A1 _07109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11207__A2 register_file\[13\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12883__I _07409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15589_ _03082_ _03086_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_13_clk clknet_5_2__leaf_clk clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08130_ _03461_ _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08084__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16579__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10966__A1 _06203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08061_ _03392_ _03225_ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07831__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10718__A1 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09584__A1 _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08387__A2 _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13380__A2 _07718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10194__A2 register_file\[21\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08601__I _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08963_ _04149_ register_file\[7\]\[5\] _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09336__A1 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13132__A2 _07568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07914_ _03247_ _01010_ _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08894_ _04149_ register_file\[15\]\[4\] _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11143__A1 _06156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15409__A1 _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07845_ _03159_ _03178_ _03179_ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11694__A2 _06656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12891__A1 _07414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15434__I _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07776_ _03027_ register_file\[13\]\[23\] _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14632__A2 register_file\[24\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09515_ _04827_ _04828_ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11446__A2 _06506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08311__A2 _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09446_ _04759_ _04760_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09588__B _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09377_ _04690_ _04692_ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ _01455_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12946__A2 _07446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08075__A1 _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10957__A1 _06196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15946__CLK clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08259_ _03282_ register_file\[6\]\[29\] _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_137_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11270_ _06072_ _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10709__A1 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09575__A1 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10221_ _05522_ _05523_ _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11382__A1 _06469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09607__I _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output78_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10152_ _05451_ _05455_ _03943_ _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08511__I _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15112__A3 _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09327__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13129__I _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10083_ _05254_ register_file\[24\]\[22\] _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14960_ _02462_ _02463_ _02465_ _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11134__A1 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13911_ _01247_ register_file\[11\]\[3\] _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07889__A1 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14891_ _01042_ _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11872__I _06777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08667__B _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13842_ _01360_ _01271_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16561_ _00949_ clknet_leaf_165_clk register_file\[29\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13773_ _01009_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12634__A1 _07242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10985_ _06215_ _06216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15512_ _03010_ register_file\[31\]\[22\] _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12724_ _07314_ register_file\[20\]\[0\] _07315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16492_ _00880_ clknet_5_24__leaf_clk register_file\[15\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15443_ _02941_ _02609_ _02942_ _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12655_ _07264_ _07260_ _07265_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12937__A2 register_file\[18\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11606_ _06388_ _06602_ _06605_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15374_ _02869_ _02874_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12586_ _07016_ _07215_ _07218_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10948__A1 _06100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09802__A2 _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10437__B _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14325_ _01833_ _01837_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12208__I _06962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11537_ _06558_ register_file\[11\]\[12\] _06564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14256_ _01684_ register_file\[10\]\[7\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11468_ _06410_ _06520_ _06522_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13207_ _07612_ register_file\[15\]\[21\] _07617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10951__I _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10419_ _05717_ _05718_ _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14187_ _01158_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11373__A1 _06462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11399_ _06476_ register_file\[26\]\[21\] _06481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16101__CLK clknet_leaf_54_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13138_ _07572_ _07568_ _07573_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13114__A2 register_file\[16\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13069_ _07514_ register_file\[16\]\[7\] _07525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11125__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_2_clk clknet_5_0__leaf_clk clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09869__A2 _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14862__A2 _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11676__A2 _06641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12873__A1 _07359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16251__CLK clknet_leaf_269_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09300_ _04615_ _04616_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10100__A2 register_file\[20\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09231_ _04547_ _04548_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14378__A1 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15969__CLK clknet_leaf_314_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13502__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12928__A2 register_file\[18\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09162_ _04416_ register_file\[24\]\[8\] _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08057__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08113_ register_file\[7\]\[27\] _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07804__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09093_ _03879_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11022__I _06220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08044_ _03372_ _03375_ _03376_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_190_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09557__A1 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15429__I _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11364__A1 _06386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09995_ _05298_ _05301_ _04900_ _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09309__A1 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14302__A1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08780__A2 _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09871__B _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _04266_ _04267_ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14853__A2 register_file\[13\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08877_ _04198_ _04199_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11692__I _06059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15164__I _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16200__D _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07828_ _01114_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12616__A1 _07235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08296__A1 _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12092__A2 _06866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10770_ net40 _06058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09429_ _04726_ _04743_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12919__A2 _07425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12440_ _07030_ _07126_ _07130_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08048__A1 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09796__A1 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12371_ _07089_ _07090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08950__B _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14110_ _01625_ _01456_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11322_ _06383_ _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15090_ _02593_ register_file\[23\]\[17\] _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09548__A1 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13344__A2 _07697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14041_ _01018_ _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10771__I _06058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14243__I _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11253_ _06370_ _06383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_106_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11355__A1 _06454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10204_ _03831_ _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08220__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11184_ _06078_ _06337_ _06339_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16274__CLK clknet_leaf_158_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10135_ _05303_ register_file\[2\]\[22\] _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08771__A2 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15992_ _00380_ clknet_leaf_244_clk register_file\[7\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11107__A1 _06290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14943_ _02438_ _02448_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10066_ _05368_ _05371_ _05037_ _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12698__I _07247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12855__A1 _07388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11658__A2 _06630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09720__A1 _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14874_ register_file\[3\]\[14\] _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13825_ _01134_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14072__A3 _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16544_ _00932_ clknet_leaf_5_clk register_file\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13756_ _01275_ _01173_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13280__A1 _07660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12083__A2 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10968_ _06177_ _06206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12707_ _06151_ _07302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16475_ _00863_ clknet_leaf_285_clk register_file\[16\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14418__I _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11830__A2 _06751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13687_ _01206_ _01011_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10899_ _06162_ _06163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13322__I _07681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15021__A2 register_file\[13\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15426_ _02917_ _02925_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08039__A1 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12638_ _07252_ _07248_ _07253_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09021__B _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13032__A1 _07302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10167__B _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09787__A1 _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15357_ _02857_ register_file\[14\]\[20\] _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12569_ _07205_ register_file\[22\]\[15\] _07209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_5_2__f_clk_I clknet_3_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14308_ _01819_ _01475_ _01820_ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15288_ _02789_ _02542_ _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15249__I _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11777__I _06719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14239_ _01411_ register_file\[21\]\[7\] _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10149__A2 register_file\[30\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ _03771_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09780_ _04415_ _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14835__A2 register_file\[22\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15641__CLK clknet_leaf_199_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ _04053_ _04055_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12846__A1 _07276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08662_ _03889_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14599__A1 _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13941__B _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08593_ _03919_ _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15791__CLK clknet_leaf_127_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13271__A1 _07541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12074__A2 _06895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10085__A1 _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10856__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14328__I _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11821__A2 register_file\[7\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15012__A2 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13232__I _07630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09214_ _04327_ register_file\[20\]\[9\] _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16147__CLK clknet_leaf_151_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13023__A1 _07293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09145_ _04462_ _04463_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14771__A1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10388__A2 _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09076_ _04394_ _04395_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08450__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16297__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14523__A1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08027_ _03274_ register_file\[14\]\[26\] _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13326__A2 _07680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11888__A2 _06785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15079__A2 register_file\[18\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09950__A1 _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08996__I _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09978_ _05084_ register_file\[7\]\[20\] _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_301_clk_I clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14826__A2 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08929_ _03958_ register_file\[15\]\[5\] _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12837__A1 _07266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13407__I _07729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09702__A1 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12311__I _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11940_ _06818_ register_file\[5\]\[0\] _06819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10312__A2 _05613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11871_ _06769_ _06777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14054__A3 _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13610_ _01130_ register_file\[12\]\[0\] _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10822_ _06087_ register_file\[30\]\[16\] _06101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08269__A1 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13262__A1 _07531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14590_ _02099_ _01855_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12065__A2 _06888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10076__A1 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13541_ _01004_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10753_ net37 _06044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10766__I _06054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16260_ _00648_ clknet_leaf_75_clk register_file\[22\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13014__A1 _07283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13472_ _00992_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10684_ _05976_ _05979_ _03817_ _05980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15211_ register_file\[3\]\[18\] _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12423_ _07116_ register_file\[24\]\[21\] _07121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09769__A1 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16191_ _00579_ clknet_leaf_11_clk register_file\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11576__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15142_ _02644_ _01292_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12354_ _07023_ _07078_ _07079_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08441__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10715__B _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11305_ _06383_ _06420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13317__A2 _07680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15073_ _02576_ register_file\[17\]\[17\] _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08992__A2 register_file\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12285_ _06960_ register_file\[31\]\[31\] _07037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09067__I _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15664__CLK clknet_leaf_173_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14024_ register_file\[3\]\[4\] _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11236_ _06370_ _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_45_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10000__A1 _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__I _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11167_ _06321_ _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_121_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14817__A2 register_file\[31\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10118_ _03765_ _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11098_ _06283_ register_file\[27\]\[10\] _06287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15975_ _00363_ clknet_leaf_297_clk register_file\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15490__A2 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12221__I _06081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10049_ _05351_ _05354_ _04045_ _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14926_ _02430_ _02431_ _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11500__A1 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14857_ _02362_ _02112_ _02363_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15242__A2 register_file\[25\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13808_ _01096_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13253__A1 _07638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14788_ _02290_ _02295_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10067__A1 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16527_ _00915_ clknet_leaf_126_clk register_file\[14\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13739_ _01143_ register_file\[15\]\[1\] _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11803__A2 _06730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13005__A1 _07477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16458_ _00846_ clknet_5_15__leaf_clk register_file\[16\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08680__A1 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14753__A1 _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15409_ _02576_ register_file\[25\]\[21\] _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16389_ _00777_ clknet_leaf_74_clk register_file\[18\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11567__A1 _06429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_293_clk clknet_5_5__leaf_clk clknet_leaf_293_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07786__A3 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13308__A2 _07634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11319__A1 _06427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10790__A2 register_file\[30\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09901_ _05207_ _05208_ _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09832_ _04939_ register_file\[11\]\[18\] _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09763_ _04937_ register_file\[22\]\[17\] _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12819__A1 _07366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10360__B _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12131__I _06913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08714_ _03965_ register_file\[13\]\[2\] _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09694_ _05004_ register_file\[28\]\[16\] _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12295__A2 _07040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08645_ _03851_ register_file\[19\]\[1\] _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15233__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12047__A2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08576_ _03899_ _03902_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13244__A1 _07513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10058__A1 _05358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09596__B _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11558__A1 _06419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07895__I _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15687__CLK clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09128_ _04239_ register_file\[16\]\[8\] _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10230__A1 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_284_clk clknet_5_5__leaf_clk clknet_leaf_284_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ _04170_ register_file\[26\]\[7\] _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12070_ _02870_ _06895_ _06896_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_240_clk_I clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11021_ _06082_ _06236_ _06239_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09923__A1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output60_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15472__A2 _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15760_ _00148_ clknet_leaf_173_clk register_file\[13\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_255_clk_I clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12972_ _07241_ _07456_ _07463_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12286__A2 _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14711_ _02216_ _02219_ _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11923_ _06803_ register_file\[6\]\[26\] _06808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12976__I _07465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15691_ _00079_ clknet_leaf_135_clk register_file\[28\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15224__A2 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14642_ _01986_ register_file\[29\]\[12\] _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11854_ _06716_ _06722_ _06765_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12038__A2 _06874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10805_ _06028_ _06087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14573_ _02081_ _02082_ _01919_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11785_ _06647_ _06720_ _06725_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11797__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16312_ _00700_ clknet_leaf_194_clk register_file\[21\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13524_ _01023_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10736_ _06021_ _06027_ _06030_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16243_ _00631_ clknet_leaf_181_clk register_file\[23\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13455_ _07565_ _07759_ _07765_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10667_ _03920_ register_file\[11\]\[31\] _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11549__A1 _06565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12406_ _07109_ register_file\[24\]\[14\] _07111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16174_ _00562_ clknet_leaf_143_clk register_file\[25\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12210__A2 _06976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13386_ _07576_ _07718_ _07723_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10598_ _05893_ _05894_ _05895_ _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15125_ _02628_ _02378_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_275_clk clknet_5_7__leaf_clk clknet_leaf_275_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12337_ _07006_ _07064_ _07069_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15056_ _02558_ _02559_ _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12268_ _07023_ _07024_ _07025_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_208_clk_I clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14007_ _01520_ _01523_ _01148_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08717__A2 register_file\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15527__I _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11219_ _06355_ register_file\[13\]\[26\] _06360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12199_ _06970_ register_file\[31\]\[5\] _06977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11721__A1 _06675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput90 net90 rS[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_116_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15463__A2 _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12277__A2 _07024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15958_ _00346_ clknet_leaf_239_clk register_file\[8\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10288__A1 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14909_ _02414_ _02331_ _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15889_ _00277_ clknet_leaf_171_clk register_file\[11\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15262__I _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15215__A2 register_file\[1\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08430_ _03753_ _03757_ _01394_ _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12029__A2 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13226__A1 _07576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08361_ _03688_ _01059_ _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11788__A1 _06649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08292_ _01072_ register_file\[22\]\[30\] _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08653__A1 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13529__A2 _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13510__I _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10212__A1 _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10763__A2 register_file\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11960__A1 _06830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09905__A1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13701__A2 register_file\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16335__CLK clknet_leaf_146_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09435__I _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09815_ _05122_ _05123_ _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08184__A3 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09746_ _04853_ register_file\[26\]\[17\] _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12268__A2 _07024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13465__A1 _07727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09677_ _04853_ register_file\[22\]\[16\] _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16485__CLK clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15206__A2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ _03824_ register_file\[4\]\[1\] _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13217__A1 _07619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ _03777_ _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08644__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11570_ _06431_ _06582_ _06583_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12440__A2 _07126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14717__A1 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10521_ _05818_ _05819_ _05820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10451__A1 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14516__I _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13420__I _07737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13240_ _07634_ register_file\[14\]\[2\] _07637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15390__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14193__A2 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10452_ _03850_ _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08514__I _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10203__A1 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_257_clk clknet_5_16__leaf_clk clknet_leaf_257_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08947__A2 register_file\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13171_ _07590_ register_file\[15\]\[6\] _07596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10383_ _05483_ register_file\[12\]\[26\] _05684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12122_ _06926_ register_file\[3\]\[9\] _06928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12053_ _02291_ _06881_ _06886_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09345__I _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10506__A2 register_file\[26\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11004_ _06225_ register_file\[28\]\[5\] _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_194_clk_I clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15812_ _00200_ clknet_leaf_62_clk register_file\[26\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_6_0_clk clknet_0_clk clknet_3_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_74_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09124__A2 register_file\[31\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15743_ _00131_ clknet_leaf_4_clk register_file\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12955_ _07407_ register_file\[18\]\[30\] _07452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15082__I _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11906_ _06796_ register_file\[6\]\[19\] _06798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13208__A1 _07558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08883__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15674_ _00062_ clknet_leaf_257_clk register_file\[2\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12886_ _07410_ register_file\[18\]\[1\] _07412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09080__I _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15852__CLK clknet_leaf_122_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14625_ _02045_ _02132_ _02134_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11837_ _06698_ _06751_ _06756_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_89_clk_I clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14556_ _02062_ _02065_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11768_ _06712_ _06704_ _06713_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12431__A2 _07119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_132_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10442__A1 _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10719_ _06012_ _06013_ _06014_ _06015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_13507_ _01012_ _01027_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14487_ _01997_ _01914_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11699_ _06068_ _06665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_12_clk_I clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16226_ _00614_ clknet_leaf_72_clk register_file\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13438_ _07548_ _07752_ _07755_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15381__A1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14184__A2 register_file\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12195__A1 _06972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_248_clk clknet_5_16__leaf_clk clknet_leaf_248_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08938__A2 register_file\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16157_ _00545_ clknet_leaf_35_clk register_file\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_147_clk_I clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09060__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13369_ _07708_ register_file\[29\]\[22\] _07714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13931__A2 _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11942__A1 _06818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16358__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15108_ _02608_ _02609_ _02611_ _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_16088_ _00476_ clknet_leaf_235_clk register_file\[4\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_27_clk_I clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14161__I _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15039_ _01169_ _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07930_ _03262_ _03263_ _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12498__A2 register_file\[23\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13695__A1 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09363__A2 register_file\[13\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08166__A3 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07861_ _03194_ _02945_ _03195_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09600_ _04781_ register_file\[26\]\[15\] _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11170__A2 _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13447__A1 _07756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07792_ _03122_ _03127_ _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09115__A2 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09531_ _03933_ register_file\[4\]\[14\] _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13505__I _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09462_ _04763_ _04776_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08413_ _03701_ register_file\[16\]\[31\] _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_145_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10681__A1 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09393_ _04695_ _04708_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08344_ _03380_ register_file\[2\]\[30\] _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_178_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12422__A2 _07119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10864__I _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08275_ _03603_ _03604_ _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14175__A2 register_file\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_239_clk clknet_5_20__leaf_clk clknet_leaf_239_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08929__A2 register_file\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10736__A2 _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11933__A1 _06767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11695__I _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15725__CLK clknet_leaf_136_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12489__A2 register_file\[23\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13686__A1 _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09354__A2 register_file\[28\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11161__A2 _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13438__A1 _07548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15875__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _04837_ register_file\[3\]\[16\] _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13415__I _07729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12110__A1 _06652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12740_ _07250_ _07322_ _07324_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12661__A2 register_file\[21\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12671_ _07267_ register_file\[21\]\[17\] _07277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14410_ _01751_ register_file\[20\]\[9\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11622_ _06613_ register_file\[10\]\[14\] _06615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15390_ _02889_ register_file\[16\]\[21\] _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12413__A2 register_file\[24\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13610__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14341_ _01852_ _01853_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10424__A1 _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11553_ _06414_ _06568_ _06573_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10504_ _05674_ register_file\[24\]\[28\] _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14272_ _01354_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11484_ _06531_ register_file\[12\]\[23\] _06532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07840__A2 register_file\[31\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16500__CLK clknet_leaf_174_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16011_ _00399_ clknet_leaf_250_clk register_file\[6\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13223_ _07583_ register_file\[15\]\[28\] _07626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10435_ _05668_ register_file\[11\]\[27\] _05735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10727__A2 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11924__A1 _06706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09593__A2 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13154_ _07582_ _07585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10366_ _05666_ register_file\[6\]\[26\] _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15077__I _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10723__B _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12105_ _06647_ _06912_ _06917_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13085_ _06080_ _07536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10297_ _05597_ _05598_ _05599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12036_ _01704_ _06874_ _06876_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15418__A2 register_file\[28\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13429__A1 _07538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09803__I _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12101__A1 _06638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13987_ _01496_ _01503_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15726_ _00114_ clknet_leaf_146_clk register_file\[27\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12938_ _07288_ _07439_ _07442_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12652__A2 _07260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10663__A1 _05930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14929__A1 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15657_ _00045_ clknet_leaf_94_clk register_file\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12869_ _07395_ register_file\[1\]\[27\] _07401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14608_ register_file\[7\]\[11\] _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12404__A2 register_file\[24\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15588_ _03083_ _03085_ _02751_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10415__A1 _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14156__I _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09281__A1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14539_ _01800_ register_file\[1\]\[10\] _01801_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08084__A2 register_file\[28\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13060__I _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10966__A2 register_file\[2\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16180__CLK clknet_leaf_162_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15354__A1 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14157__A2 _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08060_ _03390_ _03391_ _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07831__A2 register_file\[27\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12168__A1 _06710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16209_ _00597_ clknet_leaf_155_clk register_file\[24\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15748__CLK clknet_leaf_69_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09033__A1 _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09584__A2 register_file\[22\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08962_ _04146_ register_file\[6\]\[5\] _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13668__A1 _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09336__A2 register_file\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15898__CLK clknet_leaf_265_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07913_ _03246_ _03163_ _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08893_ _04146_ register_file\[14\]\[4\] _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15409__A2 register_file\[25\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11143__A2 _06307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07844_ _01104_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12891__A2 register_file\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07775_ _02940_ register_file\[12\]\[23\] _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10859__I _06025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13235__I _07633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09514_ _04558_ register_file\[8\]\[13\] _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13840__A1 _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09445_ _04691_ register_file\[27\]\[12\] _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14396__A2 _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09376_ _04691_ register_file\[11\]\[11\] _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15593__A1 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10406__A1 _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08327_ _01162_ register_file\[14\]\[30\] _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08075__A2 register_file\[24\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10957__A2 register_file\[2\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15345__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08258_ _03580_ _03587_ _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07822__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12159__A1 _06701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08189_ _03517_ _03519_ _03369_ _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08999__I _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11906__A1 _06796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ _05254_ register_file\[20\]\[24\] _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11382__A2 register_file\[26\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10151_ _05453_ _05454_ _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09327__A2 register_file\[24\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10082_ _05252_ register_file\[25\]\[22\] _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14320__A2 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12331__A1 _07061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11134__A2 register_file\[27\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13910_ _01425_ _01427_ _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14890_ _02230_ register_file\[27\]\[15\] _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13841_ register_file\[5\]\[2\] _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14084__A1 _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16053__CLK clknet_leaf_233_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16560_ _00948_ clknet_leaf_164_clk register_file\[29\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08838__A1 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13772_ _01290_ _01006_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12634__A2 register_file\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10984_ _06214_ _06215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15511_ _01142_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10645__A1 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12723_ _07313_ _07314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_43_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16491_ _00879_ clknet_5_24__leaf_clk register_file\[15\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12654_ _07255_ register_file\[21\]\[12\] _07265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15442_ _02610_ register_file\[13\]\[21\] _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12398__A1 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11605_ _06598_ register_file\[10\]\[7\] _06605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12585_ _07212_ register_file\[22\]\[22\] _07218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15373_ _02871_ _02873_ _02544_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_168_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10948__A2 _06192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15336__A1 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14324_ _01834_ _01836_ _01494_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11536_ _06398_ _06561_ _06563_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14139__A2 _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14255_ _01682_ register_file\[11\]\[7\] _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11467_ _06517_ register_file\[12\]\[16\] _06522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09015__A1 _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13206_ _07555_ _07615_ _07616_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10418_ _05583_ register_file\[19\]\[27\] _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14186_ _01700_ _01355_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11398_ _06419_ _06479_ _06480_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12570__A1 _06999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13137_ _07563_ register_file\[16\]\[27\] _07573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12224__I _06085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10349_ _05648_ _05649_ _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14311__A2 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13068_ _06058_ _07524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11125__A2 _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12322__A1 _06992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12019_ _06865_ _06866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14075__A1 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08829__A1 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14595__B _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16546__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15709_ _00097_ clknet_leaf_32_clk register_file\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09230_ _04416_ register_file\[16\]\[9\] _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15575__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12389__A1 _07094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09161_ _04413_ register_file\[25\]\[8\] _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08112_ _03282_ register_file\[6\]\[27\] _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__15327__A1 _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11061__A1 _06156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09092_ _04406_ _04411_ _04201_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08043_ _01034_ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14614__I register_file\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12561__A1 _07198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11364__A2 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09994_ _05299_ _05300_ _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09309__A2 register_file\[10\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08945_ _04125_ register_file\[28\]\[5\] _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12313__A1 _06982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15445__I _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08876_ _04054_ register_file\[11\]\[4\] _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input22_I new_value[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07827_ _03160_ _03161_ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14066__A1 _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14605__A3 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15913__CLK clknet_leaf_111_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09428_ _04735_ _04742_ _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15566__A1 _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09359_ _04077_ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08048__A2 register_file\[2\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11052__A1 _06254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15318__A1 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09796__A2 register_file\[3\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12370_ _07086_ _07089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_16_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_16__f_clk clknet_3_4_0_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11321_ _06138_ _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output90_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14040_ _01382_ register_file\[27\]\[5\] _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09548__A2 register_file\[28\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11252_ _06049_ _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12552__A1 _07198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16419__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10203_ _05303_ register_file\[2\]\[23\] _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11355__A2 register_file\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12044__I _06873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11183_ _06334_ register_file\[13\]\[11\] _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08220__A2 register_file\[23\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10134_ _05435_ _05438_ _05037_ _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15991_ _00379_ clknet_leaf_235_clk register_file\[7\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11107__A2 register_file\[27\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14942_ _02441_ _02446_ _02447_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10065_ _05369_ _05370_ _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12855__A2 register_file\[1\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09353__I _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16569__CLK clknet_leaf_263_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10866__A1 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14873_ _02131_ register_file\[2\]\[14\] _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14057__A1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13824_ _01132_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10618__A1 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16543_ _00931_ clknet_leaf_4_clk register_file\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09484__A1 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10967_ _06135_ _06199_ _06205_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13755_ _01267_ _01274_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12706_ _07300_ _07296_ _07301_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15557__A1 _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16474_ _00862_ clknet_leaf_253_clk register_file\[16\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10898_ net35 _06162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13686_ _01205_ _01006_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15425_ _02920_ _02923_ _02924_ _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12637_ _07242_ register_file\[21\]\[7\] _07253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13032__A2 _07494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11043__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12568_ _07193_ _07208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15356_ _01161_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09787__A2 _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07798__A1 _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12791__A1 _07311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14307_ _01564_ register_file\[29\]\[8\] _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11519_ _06545_ _06553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12499_ _07009_ _07160_ _07166_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15287_ register_file\[5\]\[19\] _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14238_ _01751_ register_file\[20\]\[7\] _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16099__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14169_ _01122_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08211__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08588__B _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08730_ _04054_ register_file\[7\]\[2\] _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12846__A2 _07384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09263__I _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08661_ _03986_ register_file\[22\]\[1\] _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15936__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14599__A2 register_file\[13\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08592_ _03830_ _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09475__A1 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13271__A2 _07649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11282__A1 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15548__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09212__B _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09213_ _04325_ register_file\[21\]\[9\] _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13023__A2 _07487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09144_ _04327_ register_file\[20\]\[8\] _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12782__A1 _07347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09075_ _04327_ register_file\[20\]\[7\] _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08026_ _03357_ _03026_ _03358_ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12534__A1 _07186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09950__A2 register_file\[18\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09977_ _05082_ register_file\[6\]\[20\] _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07961__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08928_ _03956_ register_file\[14\]\[5\] _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12837__A2 _07377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09173__I _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09702__A2 register_file\[17\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08859_ _04180_ _04181_ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11870_ _06652_ _06768_ _06776_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10821_ _06099_ _06100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14519__I _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08269__A2 _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13262__A2 _07649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11273__A1 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13540_ _01057_ _01060_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10752_ _06041_ _06027_ _06043_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08517__I _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10268__B _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13471_ net6 _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12039__I _06865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10683_ _05977_ _05978_ _05979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13014__A2 _07487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12422_ _07011_ _07119_ _07120_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11025__A1 _06240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15210_ _02548_ register_file\[2\]\[18\] _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_187_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16190_ _00578_ clknet_leaf_33_clk register_file\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12773__A1 _07340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11576__A2 _06582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16241__CLK clknet_leaf_156_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15141_ _02643_ _02393_ _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10782__I _06067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12353_ _07075_ register_file\[25\]\[25\] _07079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11304_ _06116_ _06419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15072_ _01307_ _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15809__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12284_ _06163_ _07036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_153_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12525__A1 _07135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14023_ _01278_ register_file\[2\]\[4\] _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11235_ _06367_ _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_106_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16391__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10000__A2 register_file\[1\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11166_ _06046_ _06320_ _06328_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14203__B _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _05415_ _05420_ _05421_ _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11097_ _06278_ _06286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_110_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15974_ _00362_ clknet_leaf_309_clk register_file\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08201__B _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10839__A1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10048_ _05352_ _05353_ _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14925_ _02096_ register_file\[9\]\[15\] _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11500__A2 _06498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14856_ _02027_ register_file\[15\]\[14\] _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13807_ _01325_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09457__A1 _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13253__A2 register_file\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14787_ _02292_ _02294_ _02127_ _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11999_ _06701_ _06847_ _06853_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16526_ _00914_ clknet_leaf_125_clk register_file\[14\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10067__A2 register_file\[2\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13738_ _01093_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_177_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16457_ _00845_ clknet_leaf_104_clk register_file\[16\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09209__A1 _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13005__A2 register_file\[17\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14202__A1 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13669_ _01184_ _01189_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08680__A2 register_file\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11016__A1 _06233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15408_ _02826_ register_file\[24\]\[21\] _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16388_ _00776_ clknet_leaf_75_clk register_file\[18\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14753__A2 register_file\[22\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12764__A1 _07274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11567__A2 _06575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_29__f_clk_I clknet_3_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15339_ _02593_ register_file\[23\]\[20\] _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14505__A2 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11319__A2 register_file\[19\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12516__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09900_ _04939_ register_file\[19\]\[19\] _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09831_ _04937_ register_file\[10\]\[18\] _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13508__I _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07943__A1 _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09762_ _05070_ _05071_ _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12819__A2 register_file\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08713_ _04033_ _04036_ _04037_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09693_ _03843_ _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09696__A1 _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08644_ _03848_ register_file\[18\]\[1\] _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16114__CLK clknet_leaf_229_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08575_ _03901_ register_file\[4\]\[0\] _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13244__A2 _07632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_165_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11255__A1 _06378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14992__A2 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10088__B _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11007__A1 _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11558__A2 _06575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09127_ _04237_ register_file\[17\]\[8\] _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09058_ _04376_ _04377_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10230__A2 register_file\[8\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08009_ _03333_ _03341_ _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11020_ _06233_ register_file\[28\]\[12\] _06239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07934__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output53_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08021__B _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12971_ _07462_ register_file\[17\]\[3\] _07463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14710_ _02217_ register_file\[1\]\[12\] _02218_ _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11922_ _06703_ _06806_ _06807_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11494__A1 _06436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15690_ _00078_ clknet_leaf_100_clk register_file\[28\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10777__I _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14641_ _01818_ register_file\[28\]\[12\] _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11853_ _06719_ register_file\[7\]\[31\] _06765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13153__I _07583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10804_ _06085_ _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14572_ _01835_ register_file\[18\]\[11\] _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11784_ _06722_ register_file\[7\]\[2\] _06725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12994__A1 _07264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16311_ _00699_ clknet_5_19__leaf_clk register_file\[21\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11797__A2 register_file\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13523_ _01043_ register_file\[22\]\[0\] _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10735_ _06029_ register_file\[30\]\[0\] _06030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16242_ _00630_ clknet_leaf_156_clk register_file\[23\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15631__CLK clknet_leaf_152_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10666_ _03828_ register_file\[10\]\[31\] _05962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13454_ _07763_ register_file\[9\]\[24\] _07765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12746__A1 _07326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12405_ _06994_ _07105_ _07110_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16173_ _00561_ clknet_leaf_138_clk register_file\[25\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13385_ _07679_ register_file\[29\]\[29\] _07723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09611__A1 _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10597_ _05640_ register_file\[1\]\[29\] _05895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15124_ _02622_ _02627_ _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12336_ _07068_ register_file\[25\]\[18\] _07069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15055_ _02390_ register_file\[25\]\[17\] _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12267_ _07019_ register_file\[31\]\[25\] _07025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08178__A1 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13171__A1 _07590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14006_ _01521_ _01258_ _01522_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11218_ _06139_ _06358_ _06359_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12198_ _06975_ _06976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_155_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput80 net80 rS[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_151_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput91 net91 rS[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__13328__I _07689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11721__A2 register_file\[8\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12232__I _06975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11149_ _06315_ _06316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_96_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15957_ _00345_ clknet_leaf_221_clk register_file\[8\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09678__A1 _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15543__I register_file\[5\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14908_ _02412_ _02413_ _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11485__A1 _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15888_ _00276_ clknet_leaf_186_clk register_file\[11\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14839_ _02338_ _02345_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13226__A2 _07622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16287__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08360_ register_file\[5\]\[31\] _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11237__A1 _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14974__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12985__A1 _07254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11788__A2 _06720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16509_ _00897_ clknet_leaf_300_clk register_file\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08291_ _03618_ _01084_ _03619_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08653__A2 register_file\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09850__A1 _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_300_clk_I clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12737__A1 _07318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09602__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08405__A2 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11311__I _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10212__A2 register_file\[17\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11960__A2 register_file\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15151__A2 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08169__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07916__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09814_ _04919_ register_file\[4\]\[18\] _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15454__A3 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09745_ _05053_ _05054_ _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14662__A1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13465__A2 register_file\[9\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15453__I _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09676_ _04985_ _04986_ _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08627_ _03821_ register_file\[5\]\[1\] _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14414__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13217__A2 register_file\[15\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11228__A1 _06160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15654__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08558_ _03881_ _03884_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08489_ _03815_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10520_ _05758_ register_file\[28\]\[28\] _05819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14717__A2 register_file\[25\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12728__A1 _07314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10451_ _05750_ register_file\[6\]\[27\] _05751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15390__A2 register_file\[16\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11400__A1 _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13170_ _07518_ _07594_ _07595_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10203__A2 register_file\[2\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10382_ _05481_ register_file\[13\]\[26\] _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12121_ _06662_ _06922_ _06927_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15142__A2 _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12052_ _06885_ net15 _06886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11003_ _06228_ _06229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12900__A1 _07250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15811_ _00199_ clknet_leaf_49_clk register_file\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11891__I _06769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11467__A1 _06517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15742_ _00130_ clknet_leaf_8_clk register_file\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12954_ _07304_ _07446_ _07451_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11905_ _06686_ _06792_ _06797_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15673_ _00061_ clknet_leaf_241_clk register_file\[2\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14405__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13208__A2 _07615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_193_clk clknet_5_24__leaf_clk clknet_leaf_193_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12885_ _07230_ _07408_ _07411_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11219__A1 _06355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14624_ _02133_ _01883_ _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11836_ _06755_ register_file\[7\]\[23\] _06756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12967__A1 _07237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14555_ _02063_ _02064_ _01982_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09832__A1 _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11767_ _06640_ register_file\[8\]\[29\] _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13611__I _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13506_ _01016_ _01020_ _01026_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10442__A2 register_file\[15\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10718_ _03922_ register_file\[1\]\[31\] _06014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14486_ _01995_ _01996_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11698_ _06662_ _06656_ _06664_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12719__A1 _06216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16225_ _00613_ clknet_leaf_72_clk register_file\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13437_ _07749_ register_file\[9\]\[17\] _07755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15381__A2 register_file\[1\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10649_ _03880_ register_file\[13\]\[30\] _05946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12195__A2 _06961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16156_ _00544_ clknet_leaf_35_clk register_file\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13368_ _07558_ _07711_ _07713_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09060__A2 register_file\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15538__I _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15107_ _02610_ register_file\[13\]\[17\] _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11942__A2 register_file\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12319_ _07054_ register_file\[25\]\[11\] _07059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14442__I _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16087_ _00475_ clknet_leaf_234_clk register_file\[4\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13299_ _07667_ register_file\[14\]\[26\] _07672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13144__A1 _07576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08440__I _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15038_ _02541_ _02542_ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09899__A1 _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14892__A1 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13695__A2 register_file\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07860_ _02859_ register_file\[15\]\[24\] _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09980__B _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07791_ _03124_ _03126_ _02960_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14644__A1 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13447__A2 register_file\[9\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11458__A1 _06400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09530_ _04809_ _04843_ _04641_ net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09461_ _04770_ _04775_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08412_ _03730_ _03739_ _01468_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09392_ _04702_ _04707_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14947__A2 _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12958__A1 _07308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08343_ _03671_ _01052_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14617__I _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11630__A1 _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08274_ _03459_ register_file\[1\]\[29\] _01198_ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15372__A2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_254_clk_I clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13383__A1 _07679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16302__CLK clknet_leaf_145_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13922__A3 _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11976__I _06825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10880__I _06147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13135__A1 _07570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14883__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_269_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13686__A2 _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16452__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11697__A1 _06663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15427__A3 _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13438__A2 _07752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07989_ _03319_ _03155_ _03321_ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11449__A1 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09728_ _04967_ register_file\[2\]\[16\] _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12110__A2 _06912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_175_clk clknet_5_29__leaf_clk clknet_leaf_175_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10121__A1 _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09659_ _04970_ register_file\[1\]\[15\] _04971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11216__I _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10120__I _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12670_ _06103_ _07276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15060__A1 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_207_clk_I clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12949__A1 _07443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11621_ _06402_ _06609_ _06614_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15132__B _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09814__A1 _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11621__A1 _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14340_ _01423_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11552_ _06572_ register_file\[11\]\[18\] _06573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10276__B _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08093__A3 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10503_ _05672_ register_file\[25\]\[28\] _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14271_ register_file\[7\]\[7\] _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11483_ _06494_ _06531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13374__A1 _07715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16010_ _00398_ clknet_leaf_292_clk register_file\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13222_ _07572_ _07622_ _07625_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10434_ _05666_ register_file\[10\]\[27\] _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15358__I _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11924__A2 _06806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14262__I _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13153_ _07583_ _07584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10365_ _04316_ _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12104_ _06914_ register_file\[3\]\[2\] _06917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13084_ _07534_ _07532_ _07535_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08260__I register_file\[7\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10296_ _05397_ register_file\[8\]\[25\] _05598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12035_ _06870_ net39 _06876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11688__A1 _06654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14626__A1 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13429__A2 _07745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13986_ _01499_ _01502_ _01237_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12101__A2 _06912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15725_ _00113_ clknet_leaf_136_clk register_file\[27\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12937_ _07436_ register_file\[18\]\[22\] _07442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10112__A1 _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_166_clk clknet_5_31__leaf_clk clknet_leaf_166_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15656_ _00044_ clknet_leaf_94_clk register_file\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11860__A1 _06770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12868_ _07298_ _07398_ _07400_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15051__A1 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14607_ _02033_ register_file\[6\]\[11\] _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_21_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11819_ _06741_ register_file\[7\]\[16\] _06746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15587_ _03084_ register_file\[18\]\[23\] _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12799_ _06317_ _03927_ _07358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14538_ _02045_ _02046_ _02048_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08435__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10415__A2 register_file\[16\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14469_ _01018_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14157__A3 _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15354__A2 register_file\[13\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16208_ _00596_ clknet_leaf_154_clk register_file\[24\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13365__A1 _07708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12168__A2 _06950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16139_ _00527_ clknet_leaf_98_clk register_file\[31\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13117__A1 _07551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08792__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08961_ _04281_ _04282_ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11679__A1 _06650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07912_ _03244_ _03245_ _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08892_ _04212_ _04214_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07843_ _03170_ _03177_ _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10351__A1 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12420__I _07097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07774_ _03105_ _03109_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ _04556_ register_file\[9\]\[13\] _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_157_clk clknet_5_31__leaf_clk clknet_leaf_157_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10103__A1 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09444_ _04689_ register_file\[26\]\[12\] _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11851__A1 _06719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10875__I _06143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ _03889_ _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15593__A2 register_file\[21\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11603__A1 _06598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08345__I register_file\[3\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10406__A2 register_file\[2\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08326_ _03653_ _03436_ _03654_ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_193_clk_I clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08257_ _03583_ _03586_ _03279_ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15345__A2 register_file\[9\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13356__A1 _07546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12159__A2 _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_5_0_clk clknet_0_clk clknet_3_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_153_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_73_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08188_ _03518_ _01167_ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13108__A1 _07550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10150_ _05248_ register_file\[31\]\[23\] _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15842__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14856__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13659__A2 _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_88_clk_I clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10081_ _05382_ _05385_ _04018_ _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08535__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12331__A2 register_file\[25\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_131_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15992__CLK clknet_leaf_244_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13840_ _01162_ _01358_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_11_clk_I clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12095__A1 _06266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_148_clk clknet_5_27__leaf_clk clknet_leaf_148_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13771_ _01288_ _01289_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10983_ _03769_ net43 _06214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_146_clk_I clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15510_ _01093_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12722_ _07310_ _07313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_74_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16490_ _00878_ clknet_leaf_114_clk register_file\[15\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10645__A2 register_file\[23\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11842__A1 _06703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15441_ _02940_ register_file\[12\]\[21\] _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12653_ _06081_ _07264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15584__A2 _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12398__A2 _07105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11604_ _06386_ _06602_ _06604_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15372_ _02872_ _02542_ _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12584_ _07014_ _07215_ _07217_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14323_ _01835_ register_file\[18\]\[8\] _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11535_ _06558_ register_file\[11\]\[11\] _06563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16498__CLK clknet_leaf_175_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15336__A2 register_file\[21\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14254_ _01767_ _01427_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11466_ _06407_ _06520_ _06521_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09015__A2 register_file\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15088__I _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13898__A2 _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13205_ _07612_ register_file\[15\]\[20\] _07616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10417_ _05452_ register_file\[18\]\[27\] _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11397_ _06476_ register_file\[26\]\[20\] _06480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14185_ register_file\[7\]\[6\] _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12570__A2 _07208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13136_ _06146_ _07572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10348_ _05449_ register_file\[16\]\[26\] _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10581__A1 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14720__I _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13067_ _07522_ _07520_ _07523_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10279_ _05579_ _05580_ _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12322__A2 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12018_ _06862_ _06865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15272__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14075__A2 register_file\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_139_clk clknet_5_26__leaf_clk clknet_leaf_139_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08829__A2 register_file\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13969_ _01308_ register_file\[17\]\[4\] _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15708_ _00096_ clknet_leaf_36_clk register_file\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11833__A1 _06748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14167__I _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15639_ _00027_ clknet_leaf_212_clk register_file\[30\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15575__A2 register_file\[31\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15715__CLK clknet_leaf_54_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13071__I _06062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12389__A2 register_file\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09160_ _04475_ _04478_ _04201_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_187_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08111_ _03434_ _03442_ _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09091_ _04408_ _04410_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15327__A2 register_file\[17\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11061__A2 _06257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13338__A1 _07694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08042_ _03373_ _03374_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15865__CLK clknet_leaf_260_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12010__A1 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12415__I _07086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12561__A2 register_file\[22\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13955__B _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09993_ _05168_ register_file\[23\]\[20\] _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10572__A1 _05854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08944_ _04122_ register_file\[29\]\[5\] _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12313__A2 _07050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10324__A1 _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08875_ _04052_ register_file\[10\]\[4\] _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07826_ _02993_ register_file\[25\]\[24\] _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15263__A1 _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14066__A2 register_file\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input15_I new_value[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13690__B _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11824__A1 _06748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ _04738_ _04741_ _04400_ _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15566__A2 register_file\[27\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13577__A1 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09358_ _04672_ _04673_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08309_ _01123_ register_file\[30\]\[30\] _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15318__A2 register_file\[29\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11052__A2 register_file\[28\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09289_ _04596_ _04605_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_302_clk clknet_5_4__leaf_clk clknet_leaf_302_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_166_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13329__A1 _07686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11320_ _06429_ _06420_ _06430_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12001__A1 _06851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11251_ _06380_ _06369_ _06381_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output83_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08756__A1 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12552__A2 register_file\[22\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10202_ _05500_ _05505_ _03992_ _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11182_ _06073_ _06337_ _06338_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10133_ _05436_ _05437_ _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15990_ _00378_ clknet_leaf_237_clk register_file\[7\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10064_ _05168_ register_file\[11\]\[21\] _05370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14941_ _01147_ _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09181__A1 _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10866__A2 _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14872_ _02377_ _02378_ _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16170__CLK clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14057__A2 register_file\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13823_ _01253_ register_file\[12\]\[2\] _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12995__I _07457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15371__I register_file\[5\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08694__B _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16542_ _00930_ clknet_leaf_302_clk register_file\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11815__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13754_ _01269_ _01272_ _01273_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10618__A2 register_file\[29\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10966_ _06203_ register_file\[2\]\[24\] _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12705_ _07291_ register_file\[21\]\[27\] _07301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16473_ _00861_ clknet_leaf_202_clk register_file\[16\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13685_ _01203_ _01204_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10897_ _06160_ _06029_ _06161_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_182_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15424_ _01670_ _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12636_ _06059_ _07252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15888__CLK clknet_leaf_186_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12240__A1 _07004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11043__A2 _06250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15355_ _02854_ _02609_ _02855_ _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12567_ _06997_ _07201_ _07207_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15309__A2 _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14306_ _01818_ register_file\[28\]\[8\] _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11518_ _06380_ _06544_ _06552_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15286_ _02786_ _02787_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12498_ _07164_ register_file\[23\]\[19\] _07166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10464__B _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12235__I _06099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14237_ _01318_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_171_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11449_ _06390_ _06506_ _06511_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08747__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14168_ _01682_ register_file\[11\]\[6\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08869__B _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13119_ _06124_ _07560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14099_ _01612_ _01614_ _01266_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15493__A1 _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16513__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input7_I addrS[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10306__A1 _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08660_ _03886_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12059__A1 _06885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08591_ _03917_ register_file\[2\]\[0\] _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_3_4_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11806__A1 _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_22__f_clk clknet_3_5_0_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08278__A3 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15548__A2 register_file\[2\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11314__I _06129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09212_ _04525_ _04528_ _04529_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14220__A2 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09143_ _04325_ register_file\[21\]\[8\] _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09074_ _04325_ register_file\[21\]\[7\] _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12782__A2 register_file\[20\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16043__CLK clknet_leaf_289_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08025_ _03027_ register_file\[13\]\[26\] _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12534__A2 register_file\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10545__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08779__B _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09976_ _05281_ _05282_ _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16193__CLK clknet_leaf_70_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07961__A2 register_file\[2\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08927_ _04247_ _04248_ _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08858_ _03958_ register_file\[31\]\[4\] _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14039__A2 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08910__A1 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07809_ _03143_ _02978_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08789_ _03967_ register_file\[8\]\[3\] _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10820_ _06098_ _06099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09403__B _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12470__A1 _06980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11273__A2 _06396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10751_ _06042_ register_file\[30\]\[3\] _06043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15539__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13470_ _07580_ _07730_ _07773_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10682_ _03811_ register_file\[31\]\[31\] _05978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12421_ _07116_ register_file\[24\]\[20\] _07120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12222__A1 _06983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11025__A2 register_file\[28\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12773__A2 register_file\[20\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15140_ _02641_ _02642_ _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12352_ _07049_ _07078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_127_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10784__A1 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10284__B _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11303_ _06417_ _06408_ _06418_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15071_ _02411_ register_file\[16\]\[17\] _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12283_ _07034_ _06963_ _07035_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12525__A2 register_file\[23\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14022_ _01537_ _01538_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16536__CLK clknet_leaf_241_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11234_ _06368_ _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10536__A1 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15366__I register_file\[7\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11165_ _06326_ register_file\[13\]\[4\] _06328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15475__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14278__A2 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10116_ _03913_ _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11096_ _06069_ _06279_ _06285_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15973_ _00361_ clknet_leaf_313_clk register_file\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10047_ _05084_ register_file\[15\]\[21\] _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14924_ _02349_ register_file\[8\]\[15\] _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10839__A2 _06096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15227__A1 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08901__A1 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14855_ _02025_ register_file\[14\]\[14\] _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13614__I _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13806_ _01092_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14786_ _02293_ _02125_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09457__A2 register_file\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11998_ _06851_ register_file\[5\]\[24\] _06853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14450__A2 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16525_ _00913_ clknet_leaf_125_clk register_file\[14\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13737_ _01139_ register_file\[14\]\[1\] _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10949_ _06189_ register_file\[2\]\[17\] _06195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12461__A1 _07142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_70_clk clknet_5_10__leaf_clk clknet_leaf_70_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16456_ _00844_ clknet_leaf_86_clk register_file\[16\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09209__A2 register_file\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13668_ _01186_ register_file\[1\]\[0\] _01188_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_176_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15407_ _02898_ _02906_ _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16066__CLK clknet_leaf_310_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12213__A1 _06985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11016__A2 register_file\[28\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12619_ _07235_ register_file\[21\]\[2\] _07240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16387_ _00775_ clknet_leaf_60_clk register_file\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14445__I register_file\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13599_ _01119_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08968__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12764__A2 _07336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15338_ _02590_ register_file\[22\]\[20\] _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15269_ _02520_ register_file\[10\]\[19\] _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12516__A2 _07174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10527__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08196__A2 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09830_ _05137_ _05138_ _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15903__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07943__A2 register_file\[15\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09761_ _05004_ register_file\[20\]\[17\] _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08712_ _03894_ _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09692_ _05002_ register_file\[29\]\[16\] _05003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15218__A1 _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09696__A2 register_file\[30\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08643_ _03966_ _03968_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13524__I _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08574_ _03900_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09448__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12452__A1 _07138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16409__CLK clknet_leaf_263_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_61_clk clknet_5_8__leaf_clk clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11007__A2 _06229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10883__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08959__A1 _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09126_ _04440_ _04444_ _03943_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16559__CLK clknet_leaf_150_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09057_ _04239_ register_file\[24\]\[7\] _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ _03336_ _03339_ _03340_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09384__A1 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11191__A1 _06091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09959_ _04998_ register_file\[11\]\[20\] _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09136__A1 _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12970_ _07457_ _07462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output46_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11921_ _06803_ register_file\[6\]\[25\] _06807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11494__A2 _06534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14640_ _02145_ _02148_ _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08528__I _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11852_ _06714_ _06722_ _06764_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14432__A2 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10803_ _06084_ _06085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16089__CLK clknet_leaf_248_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14571_ _01746_ register_file\[19\]\[11\] _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12443__A1 _07087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11783_ _06645_ _06720_ _06724_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_52_clk clknet_5_8__leaf_clk clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16310_ _00698_ clknet_leaf_182_clk register_file\[21\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08111__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13522_ _01042_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12994__A2 _07473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10734_ _06028_ _06029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16241_ _00629_ clknet_leaf_156_clk register_file\[23\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07870__A1 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13453_ _07562_ _07759_ _07764_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10665_ _03703_ _03763_ _05960_ _05961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14735__A3 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09359__I _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12404_ _07109_ register_file\[24\]\[13\] _07110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12746__A2 register_file\[20\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16172_ _00560_ clknet_leaf_138_clk register_file\[25\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08263__I register_file\[4\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13384_ _07574_ _07718_ _07722_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10596_ _03832_ register_file\[3\]\[29\] _05894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10757__A1 _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15123_ _02624_ _02626_ _02544_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12335_ _07038_ _07068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15054_ _02474_ register_file\[24\]\[17\] _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12266_ _06975_ _07024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13609__I _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14005_ _01143_ register_file\[15\]\[4\] _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13171__A2 register_file\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11217_ _06355_ register_file\[13\]\[25\] _06359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12197_ _06962_ _06975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput70 net70 rD[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11182__A1 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput81 net81 rS[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput92 net92 rS[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11148_ _03764_ net43 _06315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09127__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15956_ _00344_ clknet_leaf_221_clk register_file\[8\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11079_ _06270_ _06275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09678__A2 register_file\[23\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14907_ _02159_ register_file\[17\]\[15\] _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10968__I _06177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12682__A1 _07279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15887_ _00275_ clknet_leaf_186_clk register_file\[11\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11485__A2 _06527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14838_ _02341_ _02344_ _02091_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12434__A1 _07023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14769_ _02274_ _02275_ _02276_ _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43_clk clknet_5_12__leaf_clk clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_162_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12985__A2 _07466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16508_ _00896_ clknet_leaf_287_clk register_file\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08290_ _01086_ register_file\[21\]\[30\] _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11799__I _06721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10996__A1 _06037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16439_ _00827_ clknet_leaf_204_clk register_file\[17\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_192_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12737__A2 register_file\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09602__A2 register_file\[27\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09366__A1 _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08169__A2 register_file\[8\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11173__A1 _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09813_ _04917_ register_file\[5\]\[18\] _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07916__A2 register_file\[18\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11039__I _06228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09118__A1 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14111__A1 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09744_ _04919_ register_file\[24\]\[17\] _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14662__A2 register_file\[21\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09675_ _04919_ register_file\[20\]\[16\] _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08626_ _03944_ _03951_ _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12425__A1 _07116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08557_ _03883_ register_file\[8\]\[0\] _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11228__A2 _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_34_clk clknet_5_6__leaf_clk clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08488_ _03790_ _03814_ _03792_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_35_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16381__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07852__A1 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15949__CLK clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10450_ _03847_ _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_178_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09109_ _04427_ _04428_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10118__I _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11400__A2 _06479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10381_ _05662_ _05681_ _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12120_ _06926_ register_file\[3\]\[8\] _06927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09357__A1 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14350__A1 _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12051_ _06865_ _06885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11164__A1 _06041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11002_ _06220_ _06228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12900__A2 _07418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10911__A1 _06033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15810_ _00198_ clknet_leaf_49_clk register_file\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14653__A2 _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15741_ _00129_ clknet_leaf_281_clk register_file\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10788__I _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12953_ _07407_ register_file\[18\]\[29\] _07451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11904_ _06796_ register_file\[6\]\[18\] _06797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15672_ _00060_ clknet_leaf_240_clk register_file\[2\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12884_ _07410_ register_file\[18\]\[0\] _07411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14405__A2 register_file\[19\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15602__A1 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14623_ register_file\[3\]\[11\] _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12416__A1 _07116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11835_ _06718_ _06755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11219__A2 register_file\[13\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14554_ _01980_ register_file\[26\]\[11\] _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12967__A2 _07456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11766_ _06155_ _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10978__A1 _06156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13505_ _01025_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07843__A1 _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10717_ _03832_ register_file\[3\]\[31\] _06013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14485_ _01741_ register_file\[17\]\[10\] _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11697_ _06663_ register_file\[8\]\[8\] _06664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09089__I _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12719__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16224_ _00612_ clknet_leaf_23_clk register_file\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13916__A1 _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13436_ _07546_ _07752_ _07754_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10648_ _05937_ _05944_ _05945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16155_ _00543_ clknet_leaf_39_clk register_file\[31\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10028__I _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13367_ _07708_ register_file\[29\]\[21\] _07713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10579_ _05873_ _05876_ _04191_ _05877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15106_ _01047_ _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12318_ _06987_ _07057_ _07058_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16086_ _00474_ clknet_leaf_234_clk register_file\[4\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13298_ _07567_ _07670_ _07671_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10472__B _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09348__A1 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15037_ _01166_ _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13144__A2 _07568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12249_ _06975_ _07012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09038__B _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09899__A2 register_file\[18\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08020__A1 _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10902__A1 _06164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07790_ _03125_ _02958_ _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14644__A2 register_file\[30\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12655__A1 _07264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11458__A2 _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15939_ _00327_ clknet_leaf_14_clk register_file\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09460_ _04774_ _04637_ _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08411_ _03734_ _03738_ _01022_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12407__A1 _06997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09391_ _04706_ _04637_ _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_clk clknet_5_2__leaf_clk clknet_leaf_16_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08087__A1 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08342_ _03665_ _03670_ _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12958__A2 _07410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13080__A1 _07527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10647__B _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10969__A1 _06203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14119__B _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08273_ _03294_ _03600_ _03602_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11630__A2 _06616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11322__I _06383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_13__f_clk_I clknet_3_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13383__A2 register_file\[29\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11394__A1 _06476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14332__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13135__A2 _07568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11146__A1 _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14883__A2 register_file\[24\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08011__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11697__A2 register_file\[8\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12894__A1 _07244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15464__I _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08787__B _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07988_ _03320_ register_file\[23\]\[26\] _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15621__CLK clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14635__A2 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09727_ _05033_ _05036_ _05037_ _05038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11449__A2 _06506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09658_ _03776_ _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10121__A2 register_file\[12\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14399__A1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08609_ _03935_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_103_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09589_ _04630_ register_file\[2\]\[14\] _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15771__CLK clknet_leaf_283_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11620_ _06613_ register_file\[10\]\[13\] _06614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09814__A2 register_file\[4\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12328__I _07049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07825__A1 _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11551_ _06542_ _06572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11621__A2 _06609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _05797_ _05800_ _04655_ _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14270_ _01611_ register_file\[6\]\[7\] _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_10_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16127__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11482_ _06424_ _06527_ _06530_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_195_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13221_ _07619_ register_file\[15\]\[27\] _07625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14571__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14543__I _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13374__A2 register_file\[29\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10433_ _05730_ _05732_ _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11385__A1 _06469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08541__I _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13152_ _07582_ _07583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10364_ _05663_ _05664_ _05665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12103_ _06645_ _06912_ _06916_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14323__A1 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12063__I _06862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13083_ _07527_ register_file\[16\]\[11\] _07535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10295_ _05395_ register_file\[9\]\[25\] _05597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11137__A1 _06144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08002__A1 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12034_ _01616_ _06874_ _06875_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11688__A2 _06656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12885__A1 _07230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14626__A2 register_file\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12637__A1 _07242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13985_ _01500_ _01326_ _01501_ _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09502__A1 _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_5_3__f_clk clknet_3_0_0_clk clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12936_ _07286_ _07439_ _07441_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15724_ _00112_ clknet_5_26__leaf_clk register_file\[27\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10112__A2 register_file\[6\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_314_clk_I clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15655_ _00043_ clknet_leaf_88_clk register_file\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12867_ _07395_ register_file\[1\]\[26\] _07400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13622__I _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14606_ _02106_ _02115_ _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11818_ _06679_ _06744_ _06745_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15586_ _01404_ _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12798_ _07308_ _07314_ _07357_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14537_ _02047_ _01883_ _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07816__A1 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12238__I _06103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11749_ _06698_ _06692_ _06700_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14468_ _01813_ register_file\[27\]\[10\] _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15549__I register_file\[3\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16207_ _00595_ clknet_leaf_143_clk register_file\[24\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14562__A1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13365__A2 register_file\[29\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13419_ _07529_ _07738_ _07744_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14399_ _01572_ register_file\[16\]\[9\] _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11376__A1 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16138_ _00526_ clknet_leaf_93_clk register_file\[31\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08451__I _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13117__A2 register_file\[16\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16069_ _00457_ clknet_leaf_310_clk register_file\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08960_ _04213_ register_file\[4\]\[5\] _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5_clk clknet_5_0__leaf_clk clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15644__CLK clknet_leaf_282_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07911_ _02993_ register_file\[17\]\[25\] _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11679__A2 register_file\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08891_ _04213_ register_file\[12\]\[4\] _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12876__A1 _07306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15284__I _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07842_ _03173_ _03176_ _02924_ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12701__I _06143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09512_ _04818_ _04825_ _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14093__A3 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10103__A2 register_file\[23\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11300__A1 _06414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09443_ _04755_ _04757_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15042__A2 _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09374_ _04689_ register_file\[10\]\[11\] _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08325_ _01048_ register_file\[13\]\[30\] _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12148__I _06921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08256_ _03584_ _03361_ _03585_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13356__A2 _07704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14553__A1 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14363__I register_file\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08187_ register_file\[7\]\[28\] _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13108__A2 _07544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11119__A1 _06297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10080_ _05383_ _05384_ _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12867__A1 _07395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12611__I _07231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10342__A2 _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12619__A1 _07235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13770_ _01000_ register_file\[17\]\[2\] _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13292__A1 _07667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12095__A2 _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10982_ _06164_ _06170_ _06213_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09920__I _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13831__A3 _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12721_ _07311_ _07312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_43_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11842__A2 _06758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15440_ _01018_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12652_ _07262_ _07260_ _07263_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11603_ _06598_ register_file\[10\]\[6\] _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15371_ register_file\[5\]\[20\] _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13595__A2 _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12583_ _07212_ register_file\[22\]\[21\] _07217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14322_ _01404_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11534_ _06395_ _06561_ _06562_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14253_ _01766_ _01424_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11465_ _06517_ register_file\[12\]\[15\] _06521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11358__A1 _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13204_ _07593_ _07615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_87_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15667__CLK clknet_leaf_210_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08271__I register_file\[3\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _05714_ _05715_ _05716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08223__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14184_ _01611_ register_file\[6\]\[6\] _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11396_ _06457_ _06479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13135_ _07570_ _07568_ _07571_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10347_ _05447_ register_file\[17\]\[26\] _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14847__A2 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10581__A2 register_file\[20\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13066_ _07514_ register_file\[16\]\[6\] _07523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12858__A1 _07288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10278_ _05449_ register_file\[16\]\[25\] _05580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09723__A1 _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12017_ _06863_ _06864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11530__A1 _06558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13283__A1 _07553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12086__A2 _06902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_253_clk_I clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13968_ _01056_ register_file\[16\]\[4\] _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15053__B _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15707_ _00095_ clknet_leaf_271_clk register_file\[28\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12919_ _07269_ _07425_ _07431_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11833__A2 register_file\[7\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13899_ _01413_ _01416_ _01237_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13352__I _07689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15638_ _00026_ clknet_leaf_212_clk register_file\[30\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08446__I _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13035__A1 _07455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15569_ _03062_ _03066_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16442__CLK clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11597__A1 _06598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08110_ _03438_ _03441_ _03279_ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_174_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09090_ _04409_ register_file\[11\]\[7\] _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13338__A2 register_file\[29\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14535__A1 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08041_ _00999_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11600__I _06601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11349__A1 _06366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_0_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16592__CLK clknet_leaf_176_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12010__A2 _06854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09992_ _05166_ register_file\[22\]\[20\] _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08943_ _04246_ _04264_ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_206_clk_I clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12849__A1 _07278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15228__B _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13527__I _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08874_ _04195_ _04196_ _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11521__A1 _06550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10324__A2 register_file\[27\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07825_ _02826_ register_file\[24\]\[24\] _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13274__A1 _07543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12077__A2 _06895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13813__A3 _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14358__I register_file\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11824__A2 register_file\[7\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09426_ _04739_ _04740_ _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13026__A1 _07295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09357_ _04602_ register_file\[31\]\[11\] _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14774__A1 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11588__A1 _06594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08308_ _03635_ _01133_ _03636_ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_166_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09288_ _04599_ _04604_ _03856_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13329__A2 register_file\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08239_ _03565_ _03568_ _03340_ _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_153_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11250_ _06378_ register_file\[19\]\[4\] _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10012__A1 _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10201_ _05502_ _05504_ _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08756__A2 register_file\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11181_ _06334_ register_file\[13\]\[10\] _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output76_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10132_ _05168_ register_file\[11\]\[22\] _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10570__B _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09705__A1 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08508__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14940_ _02443_ _02112_ _02445_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10063_ _05166_ register_file\[10\]\[21\] _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11512__A1 _06546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14977__B _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09181__A2 register_file\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14871_ _01146_ _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15254__A2 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13822_ _01337_ _01340_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13265__A1 _07646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10079__A1 _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13753_ _01169_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16541_ _00929_ clknet_leaf_301_clk register_file\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10965_ _06130_ _06199_ _06204_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11815__A2 _06737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12704_ _06147_ _07300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13017__A1 _07484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13684_ _01000_ register_file\[17\]\[1\] _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16472_ _00860_ clknet_5_19__leaf_clk register_file\[16\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10896_ _06026_ register_file\[30\]\[30\] _06161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15423_ _02921_ _02592_ _02922_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12635_ _07250_ _07248_ _07251_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11579__A1 _06543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15354_ _02610_ register_file\[13\]\[20\] _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12566_ _07205_ register_file\[22\]\[14\] _07207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12240__A2 _07000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10251__A1 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14305_ _01080_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14517__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11517_ _06550_ register_file\[11\]\[4\] _06552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07798__A3 _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15285_ register_file\[4\]\[19\] _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12497_ _07006_ _07160_ _07165_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14236_ _01745_ _01749_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11448_ _06510_ register_file\[12\]\[8\] _06511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09944__A1 _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14167_ _01681_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13740__A2 _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11379_ _06449_ _06469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11751__A1 _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13118_ _07558_ _07556_ _07559_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15048__B _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14098_ _01613_ _01355_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10480__B _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13347__I _07681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15493__A2 register_file\[24\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09046__B _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13049_ _07509_ _07505_ _07510_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07970__A3 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10306__A2 register_file\[14\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11503__A1 _06266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_192_clk_I clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15245__A2 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13256__A1 _07646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12059__A2 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08590_ _03916_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4_0_clk clknet_0_clk clknet_3_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_72_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14178__I _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11806__A2 _06737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13008__A1 _07484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15832__CLK clknet_leaf_260_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09211_ _03961_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09142_ _04457_ _04460_ _03962_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_130_clk_I clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10655__B _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14508__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_296_clk clknet_5_4__leaf_clk clknet_leaf_296_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09073_ _04389_ _04392_ _04323_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15982__CLK clknet_leaf_245_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11990__A1 _06691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_10_clk_I clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08024_ _03356_ register_file\[12\]\[26\] _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09935__A1 _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_145_clk_I clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11742__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10545__A2 register_file\[30\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16338__CLK clknet_leaf_162_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09975_ _05148_ register_file\[4\]\[20\] _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08926_ _04031_ register_file\[12\]\[5\] _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13495__A1 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08857_ _03956_ register_file\[30\]\[4\] _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16488__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08795__B _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07808_ _03142_ _02808_ _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_220_clk clknet_5_20__leaf_clk clknet_leaf_220_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08788_ _03965_ register_file\[9\]\[3\] _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11505__I _06543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10750_ _06028_ _06042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12470__A2 _07146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09409_ _04722_ _04723_ _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10481__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14816__I _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10681_ _03808_ register_file\[30\]\[31\] _05977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12420_ _07097_ _07119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_142_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08426__A1 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12222__A2 register_file\[31\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_287_clk clknet_5_5__leaf_clk clknet_leaf_287_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10233__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12351_ _07021_ _07071_ _07077_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10784__A2 register_file\[30\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11302_ _06415_ register_file\[19\]\[19\] _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11981__A1 _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15070_ _02566_ _02573_ _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12282_ _06960_ register_file\[31\]\[30\] _07035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14021_ _01146_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09926__A1 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11233_ _06367_ _06368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11164_ _06041_ _06320_ _06327_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13167__I _07585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10115_ _05417_ _05419_ _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15705__CLK clknet_leaf_199_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07952__A3 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11095_ _06283_ register_file\[27\]\[9\] _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15972_ _00360_ clknet_leaf_313_clk register_file\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14923_ _02410_ _02428_ _02347_ _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10046_ _05082_ register_file\[14\]\[21\] _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15227__A2 register_file\[18\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_211_clk clknet_5_23__leaf_clk clknet_leaf_211_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14854_ _02359_ _02192_ _02360_ _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13238__A1 _07634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15855__CLK clknet_leaf_127_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13805_ _01323_ register_file\[30\]\[2\] _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11997_ _06698_ _06847_ _06852_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14785_ register_file\[5\]\[13\] _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16524_ _00912_ clknet_leaf_123_clk register_file\[14\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10948_ _06100_ _06192_ _06194_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13736_ _01254_ _01133_ _01255_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12461__A2 register_file\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14738__A1 _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16455_ _00843_ clknet_leaf_64_clk register_file\[16\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10879_ _06146_ _06147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13667_ _01187_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13630__I _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15406_ _02901_ _02905_ _02658_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12618_ _06036_ _07239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08417__A1 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12213__A2 _06976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16386_ _00774_ clknet_leaf_60_clk register_file\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13598_ _01013_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13410__A1 _07518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08968__A2 register_file\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_278_clk clknet_5_6__leaf_clk clknet_leaf_278_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12549_ _07190_ register_file\[22\]\[7\] _07197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15337_ _02836_ _02672_ _02837_ _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09090__A1 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11150__I _06316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11972__A1 _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15163__A1 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15268_ _02518_ register_file\[11\]\[19\] _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13713__A2 _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14219_ _01564_ register_file\[29\]\[7\] _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15199_ _02450_ register_file\[6\]\[18\] _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_6_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11724__A1 _06675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09760_ _05002_ register_file\[21\]\[17\] _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08711_ _04034_ _04035_ _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09691_ _03964_ _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_202_clk clknet_5_19__leaf_clk clknet_leaf_202_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08642_ _03967_ register_file\[16\]\[1\] _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09504__B _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13229__A1 _07583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08573_ _03770_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11325__I _06143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14441__A3 _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12452__A2 register_file\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14729__A1 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08120__A3 _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13401__A1 _07511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ _04442_ _04443_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10215__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_269_clk clknet_5_7__leaf_clk clknet_leaf_269_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_194_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08959__A2 register_file\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13952__A2 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11963__A1 _06665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09056_ _04237_ register_file\[25\]\[7\] _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11995__I _06814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09908__A1 _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08007_ _01670_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14901__A1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15728__CLK clknet_leaf_166_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13704__A2 _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11715__A1 _06674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11191__A2 _06337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09958_ _04996_ register_file\[10\]\[20\] _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13468__A1 _07578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15878__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09136__A2 register_file\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08909_ _04229_ _04230_ _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15416__B _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12140__A1 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09889_ _05061_ register_file\[5\]\[19\] _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15209__A2 _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11920_ _06777_ _06806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14968__A1 _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11851_ _06719_ register_file\[7\]\[30\] _06764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11235__I _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10802_ net15 _06084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14570_ _02079_ _01832_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11782_ _06722_ register_file\[7\]\[1\] _06724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08647__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12443__A2 register_file\[24\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13521_ _01017_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10733_ _06025_ _06028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_18_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16240_ _00628_ clknet_leaf_151_clk register_file\[23\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13452_ _07763_ register_file\[9\]\[23\] _07764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10664_ _03933_ register_file\[8\]\[31\] _05960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08544__I _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07870__A2 _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12403_ _07089_ _07109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10206__A1 _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16171_ _00559_ clknet_leaf_98_clk register_file\[25\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13383_ _07679_ register_file\[29\]\[28\] _07722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10595_ _05637_ register_file\[2\]\[29\] _05893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11954__A1 _06654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10757__A2 _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12334_ _07004_ _07064_ _07067_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15145__A1 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15122_ _02625_ _02542_ _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14499__A3 _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15053_ _02511_ _02557_ _02473_ net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12265_ _06138_ _07023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09375__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14004_ _01139_ register_file\[14\]\[4\] _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11216_ _06329_ _06358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_155_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12196_ _06049_ _06974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput60 net60 rD[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11182__A2 _06337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput71 net71 rD[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_64_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput82 net82 rS[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_151_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07925__A3 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput93 net93 rS[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11147_ _06164_ _06271_ _06314_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13459__A1 _07763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09127__A2 register_file\[17\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15955_ _00343_ clknet_leaf_226_clk register_file\[8\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11078_ _06037_ _06269_ _06274_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13625__I _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14906_ _02411_ register_file\[16\]\[15\] _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10029_ _05334_ register_file\[7\]\[21\] _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12682__A2 register_file\[21\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15886_ _00274_ clknet_leaf_187_clk register_file\[11\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14837_ _02342_ _02175_ _02343_ _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16033__CLK clknet_leaf_314_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14768_ _01125_ _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12434__A2 _07126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16507_ _00895_ clknet_leaf_286_clk register_file\[15\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15061__B _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10984__I _06214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13719_ _01230_ _01238_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14699_ register_file\[5\]\[12\] _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10996__A2 _06219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16183__CLK clknet_leaf_190_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15384__A1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16438_ _00826_ clknet_leaf_204_clk register_file\[17\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07861__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13934__A2 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16369_ _00757_ clknet_leaf_160_clk register_file\[1\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09063__A1 _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11945__A1 _06647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08810__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15287__I register_file\[5\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12704__I _06147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09285__I _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09366__A2 register_file\[14\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11173__A2 register_file\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09812_ _05116_ _05120_ _03838_ _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10224__I _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09743_ _04917_ register_file\[25\]\[17\] _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12122__A1 _06926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13535__I _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09674_ _04917_ register_file\[21\]\[16\] _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13870__A1 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ _03947_ _03950_ _03796_ _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08341__A3 _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08556_ _03882_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12425__A2 register_file\[24\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16526__CLK clknet_leaf_125_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08487_ net3 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07852__A2 register_file\[11\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09108_ _04149_ register_file\[31\]\[7\] _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10380_ _05671_ _05680_ _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09039_ _04288_ register_file\[2\]\[6\] _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13689__A1 _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09357__A2 register_file\[31\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12050_ _02206_ _06881_ _06884_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14350__A2 register_file\[13\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12361__A1 _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11164__A2 _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11001_ _06046_ _06219_ _06227_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07907__A3 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10911__A2 _06168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15146__B _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16056__CLK clknet_leaf_244_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12113__A1 _06918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15740_ _00128_ clknet_leaf_283_clk register_file\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12952_ _07302_ _07446_ _07450_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11903_ _06766_ _06796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15671_ _00059_ clknet_leaf_224_clk register_file\[2\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12883_ _07409_ _07410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08983__B _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15602__A2 register_file\[9\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14622_ _02131_ register_file\[2\]\[11\] _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11834_ _06696_ _06751_ _06754_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12416__A2 register_file\[24\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14553_ _01813_ register_file\[27\]\[11\] _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11765_ _06710_ _06704_ _06711_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13180__I _07593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10978__A2 _06206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10716_ _03780_ register_file\[2\]\[31\] _06012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13504_ _01024_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14484_ _01994_ register_file\[16\]\[10\] _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11696_ _06642_ _06663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16223_ _00611_ clknet_leaf_24_clk register_file\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13435_ _07749_ register_file\[9\]\[16\] _07754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10647_ _05940_ _05943_ _03837_ _05944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11927__A1 _06767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13366_ _07555_ _07711_ _07712_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16154_ _00542_ clknet_leaf_269_clk register_file\[31\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10578_ _05874_ _05875_ _05876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15105_ _01774_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12317_ _07054_ register_file\[25\]\[10\] _07058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16085_ _00473_ clknet_leaf_233_clk register_file\[4\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13297_ _07667_ register_file\[14\]\[25\] _07671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09348__A2 register_file\[23\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12248_ _06116_ _07011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15036_ register_file\[5\]\[16\] _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14341__A2 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12179_ _06959_ _06962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10902__A2 _06029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12104__A1 _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15938_ _00326_ clknet_leaf_4_clk register_file\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12655__A2 _07260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16549__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10666__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15869_ _00257_ clknet_leaf_280_clk register_file\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15570__I _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08410_ _03735_ _03737_ _01159_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09390_ _04703_ _04704_ _04705_ _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12407__A2 _07105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08341_ _03667_ _03669_ _03376_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10418__A1 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09284__A1 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08087__A2 register_file\[30\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10969__A2 register_file\[2\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15357__A1 _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11091__A1 _06060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08272_ _03601_ _01156_ _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09036__A1 _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13907__A2 _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11918__A1 _06803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15109__A1 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14580__A2 _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10663__B _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12591__A1 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08133__B _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12343__A1 _07068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16079__CLK clknet_leaf_234_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07972__B _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08011__A2 register_file\[8\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12894__A2 _07408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input38_I new_value[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07987_ _01649_ _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14096__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09726_ _04001_ _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10657__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08314__A3 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09657_ _04837_ register_file\[3\]\[15\] _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15916__CLK clknet_leaf_122_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08608_ _03934_ _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_55_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09588_ _04896_ _04899_ _04900_ _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14399__A2 register_file\[16\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15596__A1 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08539_ _03862_ _03865_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12609__I _07231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08078__A2 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11550_ _06412_ _06568_ _06571_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11082__A1 _06275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07825__A2 register_file\[24\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10501_ _05798_ _05799_ _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14824__I _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11481_ _06524_ register_file\[12\]\[22\] _06530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11909__A1 _06796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13220_ _07570_ _07622_ _07624_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09578__A2 _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10432_ _05731_ register_file\[8\]\[27\] _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08822__I _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14045__B _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12582__A1 _07011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13151_ _06265_ _03875_ _07582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10363_ _05397_ register_file\[4\]\[26\] _05664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12102_ _06914_ register_file\[3\]\[1\] _06916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14323__A2 register_file\[18\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13082_ _06076_ _07534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10294_ _05586_ _05595_ _05596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12334__A1 _07004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11137__A2 _06307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12033_ _06870_ net38 _06875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08002__A2 register_file\[29\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12885__A2 _07408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09750__A2 _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10896__A1 _06026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10799__I _06081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13175__I _07585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12637__A2 register_file\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13984_ _01327_ register_file\[23\]\[4\] _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15723_ _00111_ clknet_leaf_136_clk register_file\[27\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10648__A1 _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12935_ _07436_ register_file\[18\]\[21\] _07441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15654_ _00042_ clknet_leaf_88_clk register_file\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15587__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12866_ _07295_ _07398_ _07399_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07901__I _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14605_ _02110_ _02114_ _02030_ _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08069__A2 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11817_ _06741_ register_file\[7\]\[15\] _06745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09266__A1 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15585_ _02998_ register_file\[19\]\[23\] _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12797_ _07311_ register_file\[20\]\[31\] _07357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11073__A1 _06271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15339__A1 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14536_ register_file\[3\]\[10\] _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11748_ _06699_ register_file\[8\]\[23\] _06700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09018__A1 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14734__I _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14467_ _01977_ _01811_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11679_ _06650_ register_file\[8\]\[3\] _06651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16206_ _00594_ clknet_leaf_143_clk register_file\[24\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13418_ _07742_ register_file\[9\]\[9\] _07744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08732__I _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14562__A2 register_file\[31\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14398_ _01899_ _01909_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12573__A1 _07205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11376__A2 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_5__f_clk_I clknet_3_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16137_ _00525_ clknet_leaf_95_clk register_file\[31\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16221__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13349_ _07538_ _07697_ _07702_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16068_ _00456_ clknet_leaf_313_clk register_file\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12325__A1 _06994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15565__I _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15019_ _01129_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07910_ _03243_ register_file\[16\]\[25\] _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08890_ _03900_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12876__A2 _07362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16371__CLK clknet_leaf_211_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07841_ _03174_ _03009_ _03175_ _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10887__A1 _06152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15939__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09511_ _04821_ _04824_ _04139_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11300__A2 _06408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09442_ _04756_ register_file\[24\]\[12\] _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09373_ _03886_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14250__A1 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08128__B _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08324_ _03356_ register_file\[12\]\[30\] _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11064__A1 _06218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10811__A1 _06087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09009__A1 _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08255_ _03276_ register_file\[15\]\[29\] _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14002__A1 _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14553__A2 register_file\[27\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08186_ _03282_ register_file\[6\]\[28\] _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12564__A1 _07205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11119__A2 register_file\[27\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12867__A2 register_file\[1\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09732__A2 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14069__A1 _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09709_ _04754_ register_file\[13\]\[16\] _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10981_ _06167_ register_file\[2\]\[31\] _06213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13292__A2 register_file\[14\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12720_ _07310_ _07311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15569__A1 _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15033__A3 _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12651_ _07255_ register_file\[21\]\[11\] _07263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09248__A1 _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11602_ _06382_ _06602_ _06603_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11055__A1 _06144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12582_ _07011_ _07215_ _07216_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09799__A2 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15370_ _02786_ _02870_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14321_ _01746_ register_file\[19\]\[8\] _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11533_ _06558_ register_file\[11\]\[10\] _06562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16244__CLK clknet_leaf_181_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11464_ _06505_ _06520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14252_ _01764_ _01765_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12555__A1 _06985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11358__A2 _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13203_ _07553_ _07608_ _07614_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10415_ _05449_ register_file\[16\]\[27\] _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11395_ _06417_ _06472_ _06478_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14183_ _01687_ _01697_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08223__A2 _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16394__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10346_ _05614_ _05646_ _05647_ net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13134_ _07563_ register_file\[16\]\[26\] _07571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12307__A1 _07046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15385__I _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12802__I _07358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13065_ _06054_ _07522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10277_ _05447_ register_file\[17\]\[25\] _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12858__A2 _07391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12016_ _06862_ _06863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09487__A1 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13967_ _01473_ _01483_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13283__A2 _07656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15706_ _00094_ clknet_leaf_267_clk register_file\[28\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12918_ _07429_ register_file\[18\]\[14\] _07431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09332__B _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08727__I _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13898_ _01414_ _01326_ _01415_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12249__I _06975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09239__A1 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15637_ _00025_ clknet_leaf_211_clk register_file\[30\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12849_ _07278_ _07384_ _07389_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13035__A2 register_file\[17\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11153__I _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15568_ _03064_ _03065_ _02814_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12794__A1 _07304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14519_ _01147_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15499_ _01119_ _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08040_ register_file\[5\]\[26\] _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08462__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14535__A2 register_file\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12546__A1 _06974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11349__A2 _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09991_ _05296_ _05297_ _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13808__I _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14838__A3 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15761__CLK clknet_leaf_173_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08942_ _04253_ _04263_ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12849__A2 _07384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08873_ _04125_ register_file\[8\]\[4\] _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11328__I _06147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07824_ _03148_ _03158_ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16117__CLK clknet_leaf_221_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09478__A1 _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13274__A2 _07656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11285__A1 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10388__B _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09425_ _04602_ register_file\[23\]\[12\] _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16267__CLK clknet_leaf_138_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13026__A2 _07494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11037__A1 _06247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09356_ _04600_ register_file\[30\]\[11\] _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12785__A1 _07347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08307_ _01135_ register_file\[29\]\[30\] _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09287_ _04601_ _04603_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08238_ _03566_ _01141_ _03567_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12537__A1 _06967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08169_ _03181_ register_file\[8\]\[28\] _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08205__A2 _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10200_ _05503_ register_file\[23\]\[23\] _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10012__A2 register_file\[23\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11180_ _06329_ _06337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_313_clk_I clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07964__A1 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10131_ _05166_ register_file\[10\]\[22\] _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12622__I _07234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output69_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09705__A2 register_file\[18\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ _05366_ _05367_ _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14870_ _02370_ _02376_ _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13821_ _01338_ _01339_ _01126_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09469__A1 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11276__A1 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16540_ _00928_ clknet_leaf_282_clk register_file\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13752_ _01270_ _01271_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10964_ _06203_ register_file\[2\]\[23\] _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15006__A3 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12703_ _07298_ _07296_ _07299_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16471_ _00859_ clknet_leaf_215_clk register_file\[16\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13017__A2 register_file\[17\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14214__A1 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13683_ _01202_ register_file\[16\]\[1\] _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10895_ _06159_ _06160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11028__A1 _06240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15422_ _02593_ register_file\[31\]\[21\] _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12634_ _07242_ register_file\[21\]\[6\] _07251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14765__A2 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15634__CLK clknet_leaf_178_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12776__A1 _07286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15353_ _02524_ register_file\[12\]\[20\] _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12565_ _06994_ _07201_ _07206_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09641__A1 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14304_ _01812_ _01816_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14517__A2 register_file\[15\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11516_ _06377_ _06544_ _06551_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15284_ _01530_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12496_ _07164_ register_file\[23\]\[18\] _07165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14235_ _01747_ _01748_ _01494_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11447_ _06497_ _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11200__A1 _06348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10003__A2 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11378_ _06400_ _06465_ _06468_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14166_ _01037_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11751__A2 register_file\[8\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13117_ _07551_ register_file\[16\]\[21\] _07559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10329_ _05565_ register_file\[28\]\[25\] _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14097_ register_file\[7\]\[5\] _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08231__B _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13048_ _07507_ register_file\[16\]\[1\] _07510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12700__A1 _07295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10987__I _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14999_ _02502_ _02257_ _02503_ _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13256__A2 register_file\[14\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08457__I _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13008__A2 register_file\[17\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09880__A1 _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11019__A1 _06078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09210_ _04526_ _04527_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14408__B _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09141_ _04458_ _04459_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14194__I _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12707__I _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09632__A1 _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09072_ _04390_ _04391_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08192__I register_file\[5\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14508__A2 register_file\[10\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12519__A1 _07135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08023_ _01018_ _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11990__A2 _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13538__I _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07946__A1 _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11742__A2 _06692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09974_ _05146_ register_file\[5\]\[20\] _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08141__B _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08925_ _04029_ register_file\[13\]\[5\] _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14692__A1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08856_ _04177_ _04178_ _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input20_I new_value[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09751__I _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07807_ _03140_ _03141_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14369__I register_file\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14444__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08787_ _04107_ _04110_ _03838_ _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11258__A1 _06378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15657__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08123__A1 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output107_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09408_ _04518_ register_file\[31\]\[12\] _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10481__A2 register_file\[17\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10680_ _05974_ _05975_ _05976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12758__A1 _07333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09339_ _03961_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09623__A1 _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09198__I _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12350_ _07075_ register_file\[25\]\[24\] _07077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11430__A1 _06498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10233__A2 register_file\[11\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11301_ _06112_ _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12281_ _06159_ _07034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15172__A2 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_252_clk_I clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13183__A1 _07598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11232_ _06266_ _03855_ _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14020_ _01529_ _01536_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08830__I _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07937__A1 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12930__A1 _07436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12352__I _07049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11163_ _06326_ register_file\[13\]\[3\] _06327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10114_ _05418_ register_file\[7\]\[22\] _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11094_ _06064_ _06279_ _06284_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15971_ _00359_ clknet_leaf_314_clk register_file\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_267_clk_I clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13486__A2 _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14922_ _02420_ _02427_ _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10045_ _05349_ _05350_ _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11497__A1 _06495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09661__I _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14853_ _02193_ register_file\[13\]\[14\] _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13238__A2 register_file\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13804_ _01089_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14784_ _01954_ _02291_ _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11996_ _06851_ register_file\[5\]\[23\] _06852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16582__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12997__A1 _07266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16523_ _00911_ clknet_leaf_124_clk register_file\[14\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13735_ _01135_ register_file\[13\]\[1\] _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10947_ _06189_ register_file\[2\]\[16\] _06194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16454_ _00842_ clknet_leaf_86_clk register_file\[16\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14738__A2 register_file\[17\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13666_ net9 _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10878_ net30 _06146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_205_clk_I clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12749__A1 _07326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15405_ _02902_ _02738_ _02904_ _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12617_ _07237_ _07233_ _07238_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16385_ _00773_ clknet_leaf_59_clk register_file\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08417__A2 register_file\[18\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13597_ _01116_ _01117_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13410__A2 _07738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15336_ _02673_ register_file\[21\]\[20\] _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11421__A1 _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12548_ _06978_ _07194_ _07196_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15163__A2 register_file\[27\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15267_ _02768_ _02687_ _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12479_ _07150_ register_file\[23\]\[11\] _07155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13174__A1 _07524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14218_ _01387_ register_file\[28\]\[7\] _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14910__A2 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15198_ _02693_ _02700_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07928__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12921__A1 _07429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11724__A2 register_file\[8\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12262__I _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14149_ _01319_ register_file\[20\]\[6\] _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14674__A1 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08710_ _03958_ register_file\[11\]\[2\] _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09690_ _04995_ _05000_ _04529_ _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08353__A1 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08641_ _03843_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14426__A1 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13229__A2 register_file\[15\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08187__I register_file\[7\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08572_ _03898_ register_file\[5\]\[0\] _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08105__A1 _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09853__A1 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08915__I _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11660__A1 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13401__A2 _07728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09124_ _04233_ register_file\[31\]\[8\] _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10215__A2 register_file\[18\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11412__A1 _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16305__CLK clknet_leaf_159_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09055_ _04371_ _04374_ _04094_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15154__A2 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13165__A1 _07590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08006_ _03337_ _03009_ _03338_ _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14901__A2 register_file\[31\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07919__A1 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12912__A1 _07262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11715__A2 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09957_ _05262_ _05263_ _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14665__A1 _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13468__A2 _07730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11479__A1 _06524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08908_ _03773_ register_file\[8\]\[5\] _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09888_ _05186_ _05195_ _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08344__A1 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12140__A2 _06936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08839_ _01534_ _03763_ _04161_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11850_ _06712_ _06758_ _06763_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15090__A1 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12979__A1 _07462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10801_ _06082_ _06074_ _06083_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11781_ _06638_ _06720_ _06723_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13520_ _01032_ _01036_ _01040_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08825__I _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11651__A1 _06627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10732_ _06026_ _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_158_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12347__I _07038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13451_ _07726_ _07763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15393__A2 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10663_ _05930_ _05959_ _03935_ net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_167_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12402_ _06992_ _07105_ _07108_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16170_ _00558_ clknet_leaf_93_clk register_file\[25\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10206__A2 register_file\[1\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10594_ _05888_ _05891_ _03961_ _05892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13382_ _07572_ _07718_ _07721_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_191_clk_I clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15121_ register_file\[5\]\[17\] _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12333_ _07061_ register_file\[25\]\[17\] _07067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15145__A2 register_file\[18\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_3_0_clk clknet_0_clk clknet_3_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13156__A1 _07586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_71_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15052_ _02533_ _02556_ _02471_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08560__I _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12264_ _07021_ _07012_ _07022_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14003_ _01518_ _01343_ _01519_ _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11215_ _06135_ _06351_ _06357_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12195_ _06972_ _06961_ _06973_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput50 net50 rD[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_116_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput61 net61 rD[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_29_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15822__CLK clknet_leaf_150_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15448__A3 _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput72 net72 rD[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_95_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput83 net83 rS[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11146_ _06268_ register_file\[27\]\[31\] _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10390__A1 _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput94 net94 rS[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__14656__A1 _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13459__A2 register_file\[9\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13906__I _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_86_clk_I clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12810__I _07361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15954_ _00342_ clknet_leaf_216_clk register_file\[8\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11077_ _06271_ register_file\[27\]\[2\] _06274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14905_ _01107_ _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10028_ _04319_ _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15885_ _00273_ clknet_leaf_121_clk register_file\[11\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_196_clk clknet_5_18__leaf_clk clknet_leaf_196_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11426__I _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15972__CLK clknet_leaf_313_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14836_ _02176_ register_file\[23\]\[14\] _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14959__A2 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11890__A1 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14767_ _02103_ register_file\[10\]\[13\] _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11979_ _06837_ register_file\[5\]\[16\] _06842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_144_clk_I clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13641__I _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16506_ _00894_ clknet_leaf_254_clk register_file\[15\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09340__B _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11642__A1 _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13718_ _01233_ _01236_ _01237_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_16_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10445__A2 _05744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16328__CLK clknet_leaf_79_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14698_ _01954_ _02206_ _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_24_clk_I clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16437_ _00825_ clknet_leaf_205_clk register_file\[17\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13649_ _01169_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15384__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16368_ _00756_ clknet_leaf_161_clk register_file\[1\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13797__B _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_159_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15319_ _02817_ _02733_ _02819_ _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11945__A2 _06816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16478__CLK clknet_leaf_305_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16299_ _00687_ clknet_leaf_138_clk register_file\[21\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08810__A2 register_file\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13147__A1 _07578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13698__A2 _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09811_ _05118_ _05119_ _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10381__A1 _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09742_ _05048_ _05051_ _04037_ _05052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12720__I _07310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09673_ _04980_ _04983_ _03796_ _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_187_clk clknet_5_25__leaf_clk clknet_leaf_187_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_54_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13870__A2 register_file\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08624_ _03948_ _03949_ _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11881__A1 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08555_ _03770_ _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13551__I _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11633__A1 _06414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08486_ _03809_ _03812_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15375__A2 _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11071__I _06267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13386__A1 _07576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09107_ _04146_ register_file\[30\]\[7\] _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_111_clk clknet_5_13__leaf_clk clknet_leaf_111_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13138__A1 _07572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15845__CLK clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09038_ _04355_ _04358_ _04220_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12361__A2 register_file\[25\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11000_ _06225_ register_file\[28\]\[4\] _06227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14638__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10372__A1 _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12630__I _07247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15995__CLK clknet_leaf_288_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output51_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13310__A1 _07580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12113__A2 register_file\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12951_ _07407_ register_file\[18\]\[28\] _07450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__A1 _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_178_clk clknet_5_29__leaf_clk clknet_leaf_178_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11246__I _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11902_ _06684_ _06792_ _06795_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15670_ _00058_ clknet_leaf_225_clk register_file\[2\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12882_ _07406_ _07409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_73_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15063__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14621_ _01277_ _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11833_ _06748_ register_file\[7\]\[22\] _06754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09817__A1 _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14810__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14552_ _02061_ _01811_ _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09160__B _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11764_ _06640_ register_file\[8\]\[28\] _06711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13503_ _01022_ _01023_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10715_ _06007_ _06010_ _05028_ _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14483_ _01055_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11695_ _06063_ _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_186_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16222_ _00610_ clknet_leaf_33_clk register_file\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13377__A1 _07715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13434_ _07543_ _07752_ _07753_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10646_ _05941_ _05942_ _05943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09045__A2 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11927__A2 register_file\[6\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16153_ _00541_ clknet_leaf_191_clk register_file\[31\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13365_ _07708_ register_file\[29\]\[20\] _07712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10577_ _05752_ register_file\[27\]\[29\] _05875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15104_ _02524_ register_file\[12\]\[17\] _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12316_ _07049_ _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_182_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16084_ _00472_ clknet_leaf_230_clk register_file\[4\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13296_ _07641_ _07670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14877__A1 _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15035_ _02371_ _02539_ _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12247_ _07009_ _07000_ _07010_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12178_ _06960_ _06961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10363__A1 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14629__A1 _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16000__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11129_ _06304_ register_file\[27\]\[23\] _06305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12104__A2 register_file\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13301__A1 _07667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_169_clk clknet_5_30__leaf_clk clknet_leaf_169_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15937_ _00325_ clknet_leaf_4_clk register_file\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11863__A1 _06645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15868_ _00256_ clknet_leaf_276_clk register_file\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15054__A1 _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16150__CLK clknet_leaf_181_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14819_ _02320_ _02325_ _02242_ _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_92_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15718__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15799_ _00187_ clknet_leaf_214_clk register_file\[19\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14801__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13371__I _07678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11615__A1 _06606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08340_ _03668_ _03374_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10418__A2 register_file\[19\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09284__A2 register_file\[18\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ register_file\[3\]\[29\] _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11091__A2 _06279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15357__A2 register_file\[14\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13368__A1 _07558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09036__A2 register_file\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11918__A2 register_file\[6\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12040__A1 _06878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08795__A1 _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12591__A2 _07215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12343__A2 register_file\[25\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_28__f_clk clknet_3_7_0_clk clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_173_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10354__A1 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12450__I _07134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07986_ _03153_ register_file\[22\]\[26\] _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15293__A1 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14096__A2 register_file\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09725_ _05034_ _05035_ _05036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10106__A1 _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_22__f_clk_I clknet_3_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09656_ _04967_ register_file\[2\]\[15\] _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11854__A1 _06716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10657__A2 register_file\[3\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08607_ _03928_ _03933_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09587_ _03991_ _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15596__A2 register_file\[23\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11606__A1 _06388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08538_ _03864_ register_file\[12\]\[0\] _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11082__A2 register_file\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15348__A2 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08469_ _03795_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10500_ _05668_ register_file\[7\]\[28\] _05799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11480_ _06422_ _06527_ _06529_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11909__A2 register_file\[6\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ _03802_ _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12625__I _06045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12582__A2 _07215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output99_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13150_ _07580_ _07507_ _07581_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10362_ _05395_ register_file\[5\]\[26\] _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16023__CLK clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12101_ _06638_ _06912_ _06915_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10145__I _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13081_ _07531_ _07532_ _07533_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14840__I _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10293_ _05591_ _05594_ _04026_ _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15520__A2 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08538__A1 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12334__A2 _07064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12032_ _06873_ _06874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13456__I _07737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16173__CLK clknet_leaf_138_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13983_ _01323_ register_file\[22\]\[4\] _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15722_ _00110_ clknet_leaf_101_clk register_file\[27\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12934_ _07283_ _07439_ _07440_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11845__A1 _06755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10648__A2 _05944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08710__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15653_ _00041_ clknet_leaf_69_clk register_file\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14287__I _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12865_ _07395_ register_file\[1\]\[25\] _07399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15587__A2 register_file\[18\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14604_ _02111_ _02112_ _02113_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11816_ _06729_ _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15584_ _03081_ _01010_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09266__A2 register_file\[20\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12796_ _07306_ _07314_ _07356_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14535_ _01713_ register_file\[2\]\[10\] _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15339__A2 register_file\[23\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12270__A1 _07019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11747_ _06639_ _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14466_ _01975_ _01976_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11678_ _06642_ _06650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_179_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14011__A2 _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16205_ _00593_ clknet_leaf_138_clk register_file\[24\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13417_ _07526_ _07738_ _07743_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12022__A1 _06866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10629_ _03908_ register_file\[19\]\[30\] _05926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14397_ _01903_ _01908_ _01825_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12573__A2 register_file\[22\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16136_ _00524_ clknet_leaf_90_clk register_file\[31\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13770__A1 _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13348_ _07701_ register_file\[29\]\[13\] _07702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10584__A1 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08241__A3 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10055__I _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14750__I _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16067_ _00455_ clknet_leaf_310_clk register_file\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13279_ _07630_ _07660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12325__A2 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15018_ _02517_ _02522_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16516__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10336__A1 _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07840_ _03010_ register_file\[31\]\[24\] _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10887__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15275__A1 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14078__A2 _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12089__A1 _06863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09510_ _04822_ _04823_ _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11836__A1 _06755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15027__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09441_ _04415_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15578__A2 _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09372_ _04686_ _04687_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15690__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14250__A2 register_file\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08323_ _03648_ _03651_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12261__A1 _07018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_314_clk clknet_5_0__leaf_clk clknet_leaf_314_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_32_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10811__A2 register_file\[30\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08254_ _03274_ register_file\[14\]\[29\] _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09009__A2 register_file\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14002__A2 register_file\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16046__CLK clknet_leaf_245_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12013__A1 _06815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08185_ _03508_ _03515_ _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08768__A1 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12564__A2 register_file\[22\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14660__I _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07991__A2 _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10327__A1 _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12180__I _06962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14069__A2 register_file\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07969_ _01193_ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09708_ _05015_ _05018_ _03856_ _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11827__A1 _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10980_ _06160_ _06170_ _06212_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09639_ _04947_ _04950_ _04057_ _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12650_ _06077_ _07262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11601_ _06598_ register_file\[10\]\[5\] _06603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11055__A2 _06257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12581_ _07212_ register_file\[22\]\[20\] _07216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_305_clk clknet_5_1__leaf_clk clknet_leaf_305_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_169_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14320_ _01831_ _01832_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11532_ _06553_ _06561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_106_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12004__A1 _06706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14251_ _01676_ register_file\[9\]\[7\] _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11463_ _06405_ _06513_ _06519_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14544__A3 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13202_ _07612_ register_file\[15\]\[19\] _07614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12555__A2 _07194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10414_ _05447_ register_file\[17\]\[27\] _05714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14182_ _01691_ _01696_ _01608_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11394_ _06476_ register_file\[26\]\[19\] _06478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13133_ _06142_ _07570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10345_ _03934_ _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12307__A2 register_file\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13064_ _07518_ _07520_ _07521_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10276_ _05547_ _05578_ _05313_ net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09184__A1 _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12015_ _03911_ _06214_ _06862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_11__f_clk clknet_3_2_0_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11818__A1 _06679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09613__B _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13966_ _01477_ _01482_ _01395_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09487__A2 register_file\[21\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15009__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14480__A2 _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12917_ _07266_ _07425_ _07430_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15705_ _00093_ clknet_leaf_199_clk register_file\[28\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12491__A1 _07157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13897_ _01327_ register_file\[31\]\[3\] _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11434__I _06497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12848_ _07388_ register_file\[1\]\[18\] _07389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15636_ _00024_ clknet_leaf_210_clk register_file\[30\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09239__A2 register_file\[29\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__16069__CLK clknet_leaf_310_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12243__A1 _07007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15567_ _02812_ register_file\[26\]\[23\] _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12779_ _07310_ _07347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09839__I _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14518_ _02026_ _01694_ _02028_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12794__A2 _07350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08743__I _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15498_ _02996_ _02912_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10494__B _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12265__I _06138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14449_ _01146_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12546__A2 _07194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13743__A1 _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10557__A1 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16119_ _00507_ clknet_leaf_239_clk register_file\[3\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15906__CLK clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _05230_ register_file\[20\]\[20\] _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14299__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08941_ _04256_ _04261_ _04262_ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13096__I _07519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08872_ _04122_ register_file\[9\]\[4\] _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15248__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07823_ _03152_ _03157_ _03075_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13824__I _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11809__A1 _06734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10669__B _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12482__A1 _06992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11344__I _06446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_91_clk clknet_5_14__leaf_clk clknet_leaf_91_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09424_ _04600_ register_file\[22\]\[12\] _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14223__A2 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12234__A1 _06999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09355_ _04668_ _04670_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14655__I _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08306_ _01130_ register_file\[28\]\[30\] _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09286_ _04602_ register_file\[19\]\[10\] _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10796__A1 _06078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12175__I _06020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08237_ _03420_ register_file\[31\]\[29\] _03567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14526__A3 _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12537__A2 _07184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13734__A1 _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08168_ _03481_ _03498_ _03179_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08205__A3 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12903__I _07409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08099_ _03350_ register_file\[11\]\[27\] _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10130_ _05433_ _05434_ _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11519__I _06545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10061_ _05230_ register_file\[8\]\[21\] _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11963__B _06832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13820_ _01249_ register_file\[10\]\[2\] _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10579__B _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13751_ _01166_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12473__A1 _06982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11276__A2 _06396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10963_ _06166_ _06203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16211__CLK clknet_leaf_157_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11254__I _06383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_82_clk clknet_5_11__leaf_clk clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12702_ _07291_ register_file\[21\]\[26\] _07299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16470_ _00858_ clknet_leaf_216_clk register_file\[16\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13682_ _00994_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10894_ _06158_ _06159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14214__A2 register_file\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15421_ _02590_ register_file\[30\]\[21\] _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11028__A2 register_file\[28\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12633_ _06055_ _07250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12776__A2 _07343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15352_ _02849_ _02852_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12564_ _07205_ register_file\[22\]\[13\] _07206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08563__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16361__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__A2 register_file\[28\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14303_ _01814_ _01815_ _01560_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11515_ _06550_ register_file\[11\]\[3\] _06551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15283_ _02782_ _02784_ _02537_ _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12495_ _07134_ _07164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14234_ _01405_ register_file\[18\]\[7\] _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11446_ _06388_ _06506_ _06509_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13909__I _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11200__A2 register_file\[13\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14165_ _01679_ _01427_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11377_ _06462_ register_file\[26\]\[12\] _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08512__B _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13116_ _06120_ _07558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10328_ _05563_ register_file\[29\]\[25\] _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14096_ _01611_ register_file\[6\]\[5\] _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12034__B _06875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09157__A1 _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14150__A1 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13047_ _06031_ _07509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10259_ _05554_ _05561_ _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12700__A2 _07296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14998_ _02258_ register_file\[21\]\[16\] _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14453__A2 _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13949_ _01464_ _01465_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_73_clk clknet_5_10__leaf_clk clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15402__A1 _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09880__A2 register_file\[24\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15080__B _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12216__A1 _06983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11019__A2 _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14475__I _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15619_ _00007_ clknet_leaf_20_clk register_file\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14756__A3 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16599_ _00987_ clknet_leaf_223_clk register_file\[9\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09140_ _04320_ register_file\[7\]\[8\] _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13964__A1 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08473__I _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09071_ _04320_ register_file\[19\]\[7\] _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12519__A2 register_file\[23\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08022_ _03349_ _03354_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09396__A1 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08199__A2 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12723__I _07313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15469__A1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09973_ _05261_ _05279_ _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10950__A1 _06104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14141__A1 _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08924_ _04236_ _04245_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08855_ _04031_ register_file\[28\]\[4\] _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10702__A1 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16234__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13554__I _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07806_ _02805_ register_file\[17\]\[24\] _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08371__A2 _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08786_ _04108_ _04109_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input13_I new_value[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12455__A1 _06965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_64_clk clknet_5_11__leaf_clk clknet_leaf_64_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08123__A2 register_file\[2\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16384__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09871__A2 _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09407_ _04516_ register_file\[30\]\[12\] _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12758__A2 register_file\[20\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09338_ _04652_ _04653_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10769__A1 _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09623__A2 register_file\[8\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09269_ _04518_ register_file\[23\]\[10\] _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11300_ _06414_ _06408_ _06416_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13707__A1 _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12280_ _07032_ _07024_ _07033_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09387__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13729__I _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14380__A1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11231_ _06020_ _06366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12633__I _06055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11194__A1 _06095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output81_I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12930__A2 register_file\[18\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11162_ _06321_ _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10941__A1 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09139__A1 _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11249__I _06045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10113_ _03850_ _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11093_ _06283_ register_file\[27\]\[8\] _06284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15970_ _00358_ clknet_leaf_314_clk register_file\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14921_ _02423_ _02426_ _02091_ _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10044_ _05148_ register_file\[12\]\[21\] _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14852_ _02107_ register_file\[12\]\[14\] _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14435__A2 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13803_ _01320_ _01084_ _01321_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_1_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12446__A1 _07036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14783_ register_file\[4\]\[13\] _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11995_ _06814_ _06851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14986__A3 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08114__A2 _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12997__A2 _07473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16522_ _00910_ clknet_leaf_110_clk register_file\[14\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13734_ _01253_ register_file\[12\]\[1\] _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10946_ _06095_ _06192_ _06193_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09862__A2 _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14509__B _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14199__A1 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16453_ _00841_ clknet_leaf_67_clk register_file\[16\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13665_ _01185_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_177_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10877_ _06144_ _06140_ _06145_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11712__I _06085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12749__A2 register_file\[20\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15404_ _02903_ register_file\[23\]\[21\] _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13946__A1 _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12616_ _07235_ register_file\[21\]\[1\] _07238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16384_ _00772_ clknet_leaf_17_clk register_file\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13596_ _01065_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15335_ _02586_ register_file\[20\]\[20\] _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12547_ _07190_ register_file\[22\]\[6\] _07196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16107__CLK clknet_leaf_193_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15266_ _02767_ _02685_ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12478_ _06987_ _07153_ _07154_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14217_ _01727_ _01730_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13174__A2 _07594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12543__I _07185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ _06366_ _06496_ _06499_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15197_ _02696_ _02699_ _02447_ _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11185__A1 _06334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_9__f_clk clknet_3_2_0_clk clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07928__A2 register_file\[8\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12921__A2 register_file\[18\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14148_ _01659_ _01662_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16257__CLK clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14079_ _01594_ _01427_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input5_I addrD[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12685__A1 _07279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09550__A1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08640_ _03965_ register_file\[17\]\[1\] _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09073__B _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08468__I _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10160__A2 _05463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12437__A1 _07123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08571_ _03897_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_46_clk clknet_5_12__leaf_clk clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09302__A1 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08105__A2 register_file\[13\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10999__A1 _06041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07864__A1 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11660__A2 _06594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09123_ _04441_ register_file\[30\]\[8\] _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11412__A2 _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09054_ _04372_ _04373_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08005_ _03010_ register_file\[31\]\[26\] _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14362__A1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11176__A1 _06334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12912__A2 _07425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11069__I _06267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10923__A1 _06174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09956_ _05063_ register_file\[8\]\[20\] _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14665__A2 register_file\[22\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08907_ _03767_ register_file\[9\]\[5\] _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12676__A1 _07278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09887_ _05189_ _05194_ _04131_ _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13284__I _07641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09541__A1 _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08344__A2 register_file\[2\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08838_ _03933_ register_file\[4\]\[4\] _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08378__I _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10151__A2 _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12428__A1 _07123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08769_ _04091_ _04092_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_37_clk clknet_5_7__leaf_clk clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__15774__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10800_ _06065_ register_file\[30\]\[12\] _06083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15090__A2 register_file\[23\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12979__A2 register_file\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11780_ _06722_ register_file\[7\]\[0\] _06723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11100__A1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10731_ _06025_ _06026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_14_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12628__I _06049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11532__I _06553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13450_ _07560_ _07759_ _07762_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10662_ _05945_ _05958_ _05959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09002__I _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12401_ _07102_ register_file\[24\]\[12\] _07108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12600__A1 _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10148__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13381_ _07715_ register_file\[29\]\[27\] _07721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10593_ _05889_ _05890_ _05891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15120_ _02371_ _02623_ _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12332_ _07002_ _07064_ _07066_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08280__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14064__B _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14353__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15051_ _02547_ _02555_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13156__A2 register_file\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12263_ _07019_ register_file\[31\]\[24\] _07022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14002_ _01344_ register_file\[13\]\[4\] _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11214_ _06355_ register_file\[13\]\[24\] _06357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12194_ _06970_ register_file\[31\]\[4\] _06973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput51 net51 rD[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput62 net62 rD[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput73 net73 rD[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11145_ _06160_ _06271_ _06313_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput84 net84 rS[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_110_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14656__A2 register_file\[19\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput95 net95 rS[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_114_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15953_ _00341_ clknet_leaf_216_clk register_file\[8\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11076_ _06033_ _06269_ _06273_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08335__A2 _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14904_ _02401_ _02409_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10027_ _05332_ register_file\[6\]\[21\] _05333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15884_ _00272_ clknet_leaf_124_clk register_file\[11\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12419__A1 _07009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14835_ _02173_ register_file\[22\]\[14\] _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11890__A2 _06785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_28_clk clknet_5_3__leaf_clk clknet_leaf_28_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08099__A1 _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09621__B _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14766_ _02101_ register_file\[11\]\[13\] _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11978_ _06679_ _06840_ _06841_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16505_ _00893_ clknet_5_17__leaf_clk register_file\[15\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12538__I _07185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10929_ _06064_ _06178_ _06183_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13717_ _01100_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11642__A2 _06623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14697_ register_file\[4\]\[12\] _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13919__A1 _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16436_ _00824_ clknet_leaf_167_clk register_file\[17\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13648_ _01033_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14592__A1 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16367_ _00755_ clknet_leaf_144_clk register_file\[1\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13579_ _01051_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_158_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15318_ _02818_ register_file\[29\]\[20\] _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16298_ _00686_ clknet_leaf_97_clk register_file\[21\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15136__A3 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14344__A1 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13147__A2 _07507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15249_ _01075_ _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11158__A1 _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15647__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10007__B _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09810_ _04913_ register_file\[23\]\[18\] _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09741_ _05049_ _05050_ _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12658__A1 _07267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08326__A2 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15797__CLK clknet_leaf_205_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09672_ _04981_ _04982_ _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08198__I register_file\[3\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11330__A1 _06436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08623_ _03811_ register_file\[27\]\[1\] _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11881__A2 _06778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_19_clk clknet_5_2__leaf_clk clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_251_clk_I clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08554_ _03880_ register_file\[9\]\[0\] _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13083__A1 _07527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07837__A1 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12830__A1 _07259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11633__A2 _06616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12448__I _07134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08485_ _03811_ register_file\[31\]\[0\] _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13386__A2 _07718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16422__CLK clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11397__A1 _06476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ _04424_ _04425_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13279__I _07630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09037_ _04356_ _04357_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12183__I _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13138__A2 _07568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12897__A1 _07414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15494__I _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08610__B _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10372__A2 register_file\[29\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_204_clk_I clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12649__A1 _07259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09939_ _05244_ _05245_ _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11527__I _06545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09514__A1 _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13310__A2 _07634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12950_ _07300_ _07446_ _07449_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10431__I _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__A2 register_file\[15\]\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output44_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11901_ _06789_ register_file\[6\]\[17\] _06795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12881_ _07407_ _07408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15063__A2 register_file\[28\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_219_clk_I clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14620_ _02129_ _01961_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11832_ _06694_ _06751_ _06753_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13074__A1 _07526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09817__A2 register_file\[7\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14810__A2 register_file\[28\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14551_ _02060_ _01976_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11763_ _06151_ _06710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12821__A1 _07366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08057__B _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13502_ net7 _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10714_ _06008_ _06009_ _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14482_ _01984_ _01992_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11694_ _06660_ _06656_ _06661_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13433_ _07749_ register_file\[9\]\[15\] _07753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16221_ _00609_ clknet_leaf_34_clk register_file\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13377__A2 register_file\[29\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10645_ _05695_ register_file\[23\]\[30\] _05942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11388__A1 _06410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16152_ _00540_ clknet_leaf_190_clk register_file\[31\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13364_ _07689_ _07711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08571__I _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15118__A3 _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10576_ _05750_ register_file\[26\]\[29\] _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12315_ _06985_ _07050_ _07056_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14326__A1 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15103_ _02603_ _02606_ _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10060__A1 _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16083_ _00471_ clknet_leaf_231_clk register_file\[4\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13295_ _07565_ _07663_ _07669_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14877__A2 register_file\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15034_ register_file\[4\]\[16\] _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12246_ _07007_ register_file\[31\]\[19\] _07010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08005__A1 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12888__A1 _07410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12177_ _06959_ _06960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11560__A1 _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10363__A2 register_file\[4\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11128_ _06267_ _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09505__A1 _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08308__A2 _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13301__A2 register_file\[14\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10341__I _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11059_ _06152_ _06257_ _06261_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15936_ _00324_ clknet_leaf_2_clk register_file\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11312__A1 _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11863__A2 _06768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15867_ _00255_ clknet_leaf_275_clk register_file\[12\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13652__I _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15054__A2 register_file\[24\]\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14818_ _02322_ _02323_ _02324_ _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15798_ _00186_ clknet_leaf_204_clk register_file\[19\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14801__A2 register_file\[24\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07819__A1 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14749_ _01132_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11615__A2 register_file\[10\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12812__A1 _07241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16445__CLK clknet_leaf_304_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08270_ _03380_ register_file\[2\]\[29\] _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_162_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13368__A2 _07711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14483__I _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16419_ _00807_ clknet_leaf_59_clk register_file\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08481__I _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12040__A2 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16595__CLK clknet_leaf_214_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10051__A1 _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09992__A1 _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8_clk clknet_5_1__leaf_clk clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_156_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14868__A2 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09744__A1 _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10354__A2 register_file\[25\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07985_ _03316_ _03150_ _03317_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11347__I _06449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09724_ _04832_ register_file\[11\]\[16\] _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15293__A2 register_file\[2\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11303__A1 _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10106__A2 _05410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13843__A3 _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09655_ _03916_ _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_83_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_190_clk_I clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11854__A2 _06722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13562__I _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08606_ _03772_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_27_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09586_ _04897_ _04898_ _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_3_2_0_clk clknet_0_clk clknet_3_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13056__A1 _07513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_70_clk_I clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08537_ _03863_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11606__A2 _06602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12178__I _06960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08468_ _03794_ _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15812__CLK clknet_leaf_62_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10290__A1 _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_85_clk_I clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08399_ register_file\[29\]\[31\] _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10430_ _05729_ register_file\[9\]\[27\] _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10042__A1 _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10361_ _05654_ _05661_ _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15962__CLK clknet_leaf_253_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11790__A1 _06652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12100_ _06914_ register_file\[3\]\[0\] _06915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13080_ _07527_ register_file\[16\]\[10\] _07533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15438__B _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10292_ _05592_ _05593_ _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12031_ _06865_ _06873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_143_clk_I clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11542__A1 _06565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16318__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_23_clk_I clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11257__I _06055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13295__A1 _07565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13982_ _01497_ _01410_ _01498_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_150_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_158_clk_I clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15721_ _00109_ clknet_leaf_94_clk register_file\[27\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12933_ _07436_ register_file\[18\]\[20\] _07440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16468__CLK clknet_leaf_167_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13472__I _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15652_ _00040_ clknet_leaf_69_clk register_file\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_clk_I clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12864_ _07369_ _07398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_146_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14603_ _02027_ register_file\[15\]\[11\] _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14795__A1 _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11815_ _06677_ _06737_ _06743_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15583_ _03080_ _02746_ _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12795_ _07311_ register_file\[20\]\[30\] _07356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14534_ _01176_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11746_ _06129_ _06698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08474__A1 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12270__A2 register_file\[31\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12816__I _07369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14465_ _01005_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11677_ _06040_ _06649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11720__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09397__I _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16204_ _00592_ clknet_leaf_98_clk register_file\[24\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13416_ _07742_ register_file\[9\]\[8\] _07743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10628_ _03905_ register_file\[18\]\[30\] _05925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14396_ _01905_ _01906_ _01907_ _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12022__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10033__A1 _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16135_ _00523_ clknet_leaf_92_clk register_file\[31\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13347_ _07681_ _07701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09974__A1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10559_ _05855_ _05856_ _05857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10584__A2 register_file\[23\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11781__A1 _06638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13278_ _07548_ _07656_ _07659_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16066_ _00454_ clknet_leaf_310_clk register_file\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12551__I _07185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12229_ _06995_ register_file\[31\]\[14\] _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15017_ _02519_ _02521_ _02276_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11533__A1 _06558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10336__A2 register_file\[2\]\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11167__I _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13286__A1 _07555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12089__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15919_ _00307_ clknet_leaf_186_clk register_file\[10\]\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ _04754_ register_file\[25\]\[12\] _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09081__B _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13038__A1 _07308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08476__I _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15578__A3 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09371_ _04416_ register_file\[8\]\[11\] _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08322_ _03649_ _03650_ _01025_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12261__A2 _07012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14538__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08253_ _03581_ _03436_ _03582_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15985__CLK clknet_leaf_229_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08217__A1 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13210__A1 _07560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08184_ _03511_ _03514_ _03279_ _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10024__A1 _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14941__I _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13761__A2 _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14710__A1 _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11524__A1 _06386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10327__A2 _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input43_I we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15266__A2 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_250_clk clknet_5_16__leaf_clk clknet_leaf_250_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13277__A1 _07653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07968_ _03293_ _03301_ _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09707_ _05016_ _05017_ _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11827__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13506__B _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07899_ _03227_ _03232_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09638_ _04948_ _04949_ _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13029__A1 _07491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09569_ _04880_ _04881_ _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11600_ _06601_ _06602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12580_ _07193_ _07215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11531_ _06393_ _06554_ _06560_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10263__A1 _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12636__I _06059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14250_ _01508_ register_file\[8\]\[7\] _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11462_ _06517_ register_file\[12\]\[14\] _06519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08208__A1 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13201__A1 _07550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12004__A2 _06854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10015__A1 _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13201_ _07550_ _07608_ _07613_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09956__A1 _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08759__A2 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10413_ _05682_ _05713_ _05647_ net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_183_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14181_ _01692_ _01694_ _01695_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13752__A2 _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11393_ _06414_ _06472_ _06477_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09945__I _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13132_ _07567_ _07568_ _07569_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16140__CLK clknet_leaf_139_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10344_ _05629_ _05645_ _05646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15708__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13063_ _07514_ register_file\[16\]\[5\] _07521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12371__I _07089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10275_ _05562_ _05577_ _05578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_191_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11515__A1 _06550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12014_ _06716_ _06818_ _06861_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09184__A2 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10105__B _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14800__B _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15257__A2 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_241_clk clknet_5_17__leaf_clk clknet_leaf_241_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13268__A1 _07653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15858__CLK clknet_leaf_171_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14298__I _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11818__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13965_ _01479_ _01480_ _01481_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15704_ _00092_ clknet_leaf_196_clk register_file\[28\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12916_ _07429_ register_file\[18\]\[13\] _07430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08695__A1 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12491__A2 register_file\[23\]\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13896_ _01323_ register_file\[30\]\[3\] _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15635_ _00023_ clknet_leaf_178_clk register_file\[30\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12847_ _07358_ _07388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13930__I register_file\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08447__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12243__A2 register_file\[31\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15566_ _03063_ register_file\[27\]\[23\] _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13440__A1 _07756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12778_ _07288_ _07343_ _07346_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14517_ _02027_ register_file\[15\]\[10\] _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11729_ _06107_ _06686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15497_ _02995_ _02746_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14448_ _01953_ _01959_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14379_ _01635_ register_file\[24\]\[9\] _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10557__A2 register_file\[9\]\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16118_ _00506_ clknet_leaf_238_clk register_file\[3\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12281__I _06159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ _03837_ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16049_ _00437_ clknet_leaf_230_clk register_file\[5\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08871_ _04176_ _04193_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14710__B _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15592__I _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07822_ _03154_ _03155_ _03156_ _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_29_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13259__A1 _07529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11809__A2 register_file\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08686__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12482__A2 _07153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09423_ _04736_ _04737_ _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14759__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14936__I _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15420__A2 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09354_ _04669_ register_file\[28\]\[11\] _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12234__A2 _07000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13431__A1 _07541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10245__A1 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08305_ _03630_ _03633_ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_299_clk clknet_5_4__leaf_clk clknet_leaf_299_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09285_ _03907_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13982__A2 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11360__I _06457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10796__A2 _06074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11993__A1 _06844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08236_ _01123_ register_file\[30\]\[29\] _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16163__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09938__A1 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08167_ _03490_ _03497_ _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11745__A1 _06696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08610__A1 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08098_ _03429_ _03104_ _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15487__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10060_ _05228_ register_file\[9\]\[21\] _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12170__A1 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_223_clk clknet_5_21__leaf_clk clknet_leaf_223_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10720__A2 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14998__A1 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10962_ _06126_ _06199_ _06202_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13750_ register_file\[5\]\[1\] _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08677__A1 _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12473__A2 _07146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12701_ _06143_ _07298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10484__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10893_ net34 _06158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13681_ _01106_ _01196_ _01201_ net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13750__I register_file\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15411__A2 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15420_ _02918_ _02672_ _02919_ _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12632_ _07246_ _07248_ _07249_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13422__A1 _07531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10236__A1 _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12563_ _07185_ _07205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15351_ _02850_ _02851_ _02691_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11270__I _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11984__A1 _06844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08065__B _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14302_ _01557_ register_file\[26\]\[8\] _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11514_ _06545_ _06550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12494_ _07004_ _07160_ _07163_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15282_ _02783_ _02620_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09929__A1 _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14581__I _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14233_ _01746_ register_file\[19\]\[7\] _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11445_ _06502_ register_file\[12\]\[7\] _06509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13725__A2 _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14164_ _01678_ _01424_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11376_ _06398_ _06465_ _06467_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15478__A2 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13115_ _07555_ _07556_ _07557_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10327_ _05621_ _05628_ _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14095_ _01151_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09157__A2 register_file\[10\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13046_ _07502_ _07505_ _07508_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14150__A2 register_file\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10258_ _05557_ _05560_ _04486_ _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12161__A1 _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_214_clk clknet_5_23__leaf_clk clknet_leaf_214_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10189_ _05359_ register_file\[14\]\[23\] _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14989__A1 _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16036__CLK clknet_leaf_314_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14997_ _02169_ register_file\[20\]\[16\] _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13948_ _01000_ register_file\[25\]\[4\] _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10475__A1 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08132__A3 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13879_ _01386_ _01396_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13660__I register_file\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15402__A2 register_file\[22\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15618_ _00006_ clknet_leaf_20_clk register_file\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12216__A2 register_file\[31\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13413__A1 _07734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16598_ _00986_ clknet_leaf_224_clk register_file\[9\]\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15549_ register_file\[3\]\[22\] _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11180__I _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11975__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09070_ _04317_ register_file\[18\]\[7\] _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08840__A1 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08021_ _03351_ _03353_ _03108_ _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13716__A2 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11727__A1 _06675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09396__A2 register_file\[17\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15469__A2 register_file\[1\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07946__A3 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09972_ _05269_ _05278_ _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10950__A2 _06192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08923_ _04241_ _04244_ _04102_ _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14141__A2 register_file\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13835__I _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12152__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_205_clk clknet_5_22__leaf_clk clknet_leaf_205_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08854_ _04029_ register_file\[29\]\[4\] _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07833__I _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10702__A2 register_file\[24\]\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07805_ _02889_ register_file\[16\]\[24\] _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08785_ _03958_ register_file\[23\]\[3\] _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12455__A2 _07136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16529__CLK clknet_leaf_172_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10466__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14666__I _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09406_ _04719_ _04720_ _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13404__A1 _07513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09337_ _04518_ register_file\[7\]\[11\] _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12186__I _06036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09084__A1 _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10769__A2 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11966__A1 _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _04516_ register_file\[22\]\[10\] _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08831__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08219_ _01072_ register_file\[22\]\[29\] _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09199_ _04516_ register_file\[26\]\[9\] _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11718__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11230_ _06164_ _06322_ _06365_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09387__A2 register_file\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14380__A2 register_file\[25\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11194__A2 _06344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11161_ _06037_ _06320_ _06325_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output74_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10941__A2 _06185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09139__A2 register_file\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10112_ _05416_ register_file\[6\]\[22\] _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14132__A2 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11092_ _06270_ _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16059__CLK clknet_leaf_288_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14920_ _02424_ _02175_ _02425_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10043_ _05146_ register_file\[13\]\[21\] _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13891__A1 _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14851_ _02354_ _02357_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08362__A3 _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13802_ _01086_ register_file\[29\]\[2\] _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12446__A2 _07090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13643__A1 _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14782_ _02287_ _02289_ _02120_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11994_ _06696_ _06847_ _06850_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16521_ _00909_ clknet_leaf_110_clk register_file\[14\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10457__A1 _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13733_ _01129_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10945_ _06189_ register_file\[2\]\[15\] _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15396__A1 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16452_ _00840_ clknet_leaf_67_clk register_file\[16\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08574__I _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13664_ _01003_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10876_ _06131_ register_file\[30\]\[26\] _06145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15403_ _01649_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_188_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12096__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12615_ _06032_ _07237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09075__A1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16383_ _00771_ clknet_leaf_15_clk register_file\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13595_ _01113_ _01115_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11957__A1 _06822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15334_ _02831_ _02834_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12546_ _06974_ _07194_ _07195_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15265_ _02765_ _02766_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12477_ _07150_ register_file\[23\]\[10\] _07154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15200__I register_file\[7\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14216_ _01728_ _01729_ _01560_ _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14371__A2 _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11428_ _06498_ register_file\[12\]\[0\] _06499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15196_ _02697_ _02529_ _02698_ _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_153_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11185__A2 register_file\[13\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12382__A1 _06972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11359_ _06449_ _06457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_119_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14147_ _01660_ _01661_ _01494_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08050__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15320__A1 _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14078_ _01593_ _01424_ _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12134__A1 _06933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13655__I _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13029_ _07491_ register_file\[17\]\[27\] _07497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08889__A1 _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12685__A2 register_file\[21\]\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09550__A2 register_file\[30\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11175__I _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08570_ _03764_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12437__A2 register_file\[24\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10448__A1 _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09302__A2 register_file\[27\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11903__I _06766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10999__A2 _06219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08484__I _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07864__A2 register_file\[6\]\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09066__A1 _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09122_ _03779_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11948__A1 _06649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15139__A1 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08813__A1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09053_ _04233_ register_file\[15\]\[7\] _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08004_ _03007_ register_file\[30\]\[26\] _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07828__I _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_16__f_clk_I clknet_3_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11176__A2 register_file\[13\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12373__A1 _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16201__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09955_ _05061_ register_file\[9\]\[20\] _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12125__A1 _06926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13565__I _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08906_ _04194_ _04228_ _03936_ net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12676__A2 _07272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09886_ _05191_ _05193_ _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13873__A1 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16351__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09541__A2 register_file\[26\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08837_ _04121_ _04160_ _03936_ net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11085__I _06278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15919__CLK clknet_leaf_186_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12428__A2 register_file\[24\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08768_ _03786_ register_file\[15\]\[3\] _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10439__A1 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08699_ _03811_ register_file\[23\]\[2\] _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11100__A2 register_file\[27\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10730_ _06024_ _04077_ _06025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09057__A1 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10661_ _05952_ _05957_ _05958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10429__I _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12400_ _06990_ _07105_ _07107_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13380_ _07570_ _07718_ _07720_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10592_ _03890_ register_file\[7\]\[29\] _05890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08804__A1 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12600__A2 _07222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10611__A1 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12331_ _07061_ register_file\[25\]\[16\] _07066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08280__A2 register_file\[16\]\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15050_ _02554_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12262_ _06134_ _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12364__A1 _07034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11213_ _06130_ _06351_ _06356_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14001_ _01253_ register_file\[12\]\[4\] _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12193_ _06045_ _06972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_155_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput52 net52 rD[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__15302__A1 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11144_ _06268_ register_file\[27\]\[30\] _06313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput63 net63 rD[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput74 net74 rD[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_62_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput85 net85 rS[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__12116__A1 _06658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput96 net96 rS[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15952_ _00340_ clknet_leaf_216_clk register_file\[8\]\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11075_ _06271_ register_file\[27\]\[1\] _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14903_ _02405_ _02408_ _02242_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10678__A1 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10026_ _04316_ _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_188_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09532__A2 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15883_ _00271_ clknet_leaf_121_clk register_file\[11\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15605__A2 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14834_ _02339_ _02257_ _02340_ _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_4684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12419__A2 _07112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09902__B _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14765_ _02271_ _02272_ _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08099__A2 register_file\[11\]\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11977_ _06837_ register_file\[5\]\[15\] _06841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11723__I _06099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16504_ _00892_ clknet_leaf_242_clk register_file\[15\]\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13716_ _01234_ _01094_ _01235_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10928_ _06182_ register_file\[2\]\[8\] _06183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14696_ _02201_ _02204_ _02120_ _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10850__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16435_ _00823_ clknet_leaf_167_clk register_file\[17\]\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09048__A1 _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13647_ _01165_ _01167_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13919__A2 register_file\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10859_ _06025_ _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16366_ _00754_ clknet_leaf_144_clk register_file\[1\]\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13578_ _01091_ _01094_ _01098_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15317_ _01038_ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16173__D _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12529_ _07183_ _07184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16224__CLK clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16297_ _00685_ clknet_leaf_97_clk register_file\[21\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15248_ _02667_ register_file\[26\]\[19\] _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12355__A1 _07075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09220__A1 _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15179_ _02349_ register_file\[8\]\[18\] _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12107__A1 _06918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14647__A3 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09740_ _04913_ register_file\[11\]\[17\] _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10802__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08479__I _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
.ends

