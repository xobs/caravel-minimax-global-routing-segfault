VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO minimax_rf
  CLASS BLOCK ;
  FOREIGN minimax_rf ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 800.000 ;
  PIN addrD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END addrD[0]
  PIN addrD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 4.000 ;
    END
  END addrD[1]
  PIN addrD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 4.000 ;
    END
  END addrD[2]
  PIN addrD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END addrD[3]
  PIN addrD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 4.000 ;
    END
  END addrD[4]
  PIN addrS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 0.000 70.000 4.000 ;
    END
  END addrS[0]
  PIN addrS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END addrS[1]
  PIN addrS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 0.000 85.680 4.000 ;
    END
  END addrS[2]
  PIN addrS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 0.000 93.520 4.000 ;
    END
  END addrS[3]
  PIN addrS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END addrS[4]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 0.000 360.080 4.000 ;
    END
  END clk
  PIN new_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 626.080 0.000 626.640 4.000 ;
    END
  END new_value[0]
  PIN new_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 704.480 0.000 705.040 4.000 ;
    END
  END new_value[10]
  PIN new_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 0.000 712.880 4.000 ;
    END
  END new_value[11]
  PIN new_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.160 0.000 720.720 4.000 ;
    END
  END new_value[12]
  PIN new_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 728.000 0.000 728.560 4.000 ;
    END
  END new_value[13]
  PIN new_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 0.000 736.400 4.000 ;
    END
  END new_value[14]
  PIN new_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 743.680 0.000 744.240 4.000 ;
    END
  END new_value[15]
  PIN new_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 751.520 0.000 752.080 4.000 ;
    END
  END new_value[16]
  PIN new_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 0.000 759.920 4.000 ;
    END
  END new_value[17]
  PIN new_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 767.200 0.000 767.760 4.000 ;
    END
  END new_value[18]
  PIN new_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 775.040 0.000 775.600 4.000 ;
    END
  END new_value[19]
  PIN new_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 0.000 634.480 4.000 ;
    END
  END new_value[1]
  PIN new_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 0.000 783.440 4.000 ;
    END
  END new_value[20]
  PIN new_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 790.720 0.000 791.280 4.000 ;
    END
  END new_value[21]
  PIN new_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 798.560 0.000 799.120 4.000 ;
    END
  END new_value[22]
  PIN new_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 806.400 0.000 806.960 4.000 ;
    END
  END new_value[23]
  PIN new_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 814.240 0.000 814.800 4.000 ;
    END
  END new_value[24]
  PIN new_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 822.080 0.000 822.640 4.000 ;
    END
  END new_value[25]
  PIN new_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 0.000 830.480 4.000 ;
    END
  END new_value[26]
  PIN new_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 837.760 0.000 838.320 4.000 ;
    END
  END new_value[27]
  PIN new_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 845.600 0.000 846.160 4.000 ;
    END
  END new_value[28]
  PIN new_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 0.000 854.000 4.000 ;
    END
  END new_value[29]
  PIN new_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 0.000 642.320 4.000 ;
    END
  END new_value[2]
  PIN new_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 0.000 861.840 4.000 ;
    END
  END new_value[30]
  PIN new_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 869.120 0.000 869.680 4.000 ;
    END
  END new_value[31]
  PIN new_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 0.000 650.160 4.000 ;
    END
  END new_value[3]
  PIN new_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 657.440 0.000 658.000 4.000 ;
    END
  END new_value[4]
  PIN new_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 0.000 665.840 4.000 ;
    END
  END new_value[5]
  PIN new_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 673.120 0.000 673.680 4.000 ;
    END
  END new_value[6]
  PIN new_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 0.000 681.520 4.000 ;
    END
  END new_value[7]
  PIN new_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 0.000 689.360 4.000 ;
    END
  END new_value[8]
  PIN new_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 0.000 697.200 4.000 ;
    END
  END new_value[9]
  PIN rD[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 0.000 375.760 4.000 ;
    END
  END rD[0]
  PIN rD[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 0.000 454.160 4.000 ;
    END
  END rD[10]
  PIN rD[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 0.000 462.000 4.000 ;
    END
  END rD[11]
  PIN rD[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 0.000 469.840 4.000 ;
    END
  END rD[12]
  PIN rD[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 0.000 477.680 4.000 ;
    END
  END rD[13]
  PIN rD[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 0.000 485.520 4.000 ;
    END
  END rD[14]
  PIN rD[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 492.800 0.000 493.360 4.000 ;
    END
  END rD[15]
  PIN rD[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 0.000 501.200 4.000 ;
    END
  END rD[16]
  PIN rD[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 0.000 509.040 4.000 ;
    END
  END rD[17]
  PIN rD[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 0.000 516.880 4.000 ;
    END
  END rD[18]
  PIN rD[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 0.000 524.720 4.000 ;
    END
  END rD[19]
  PIN rD[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 0.000 383.600 4.000 ;
    END
  END rD[1]
  PIN rD[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 0.000 532.560 4.000 ;
    END
  END rD[20]
  PIN rD[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 0.000 540.400 4.000 ;
    END
  END rD[21]
  PIN rD[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 0.000 548.240 4.000 ;
    END
  END rD[22]
  PIN rD[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 555.520 0.000 556.080 4.000 ;
    END
  END rD[23]
  PIN rD[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 563.360 0.000 563.920 4.000 ;
    END
  END rD[24]
  PIN rD[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 0.000 571.760 4.000 ;
    END
  END rD[25]
  PIN rD[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 0.000 579.600 4.000 ;
    END
  END rD[26]
  PIN rD[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 586.880 0.000 587.440 4.000 ;
    END
  END rD[27]
  PIN rD[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 0.000 595.280 4.000 ;
    END
  END rD[28]
  PIN rD[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 0.000 603.120 4.000 ;
    END
  END rD[29]
  PIN rD[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 0.000 391.440 4.000 ;
    END
  END rD[2]
  PIN rD[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 610.400 0.000 610.960 4.000 ;
    END
  END rD[30]
  PIN rD[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 0.000 618.800 4.000 ;
    END
  END rD[31]
  PIN rD[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 0.000 399.280 4.000 ;
    END
  END rD[3]
  PIN rD[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 0.000 407.120 4.000 ;
    END
  END rD[4]
  PIN rD[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 4.000 ;
    END
  END rD[5]
  PIN rD[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.240 0.000 422.800 4.000 ;
    END
  END rD[6]
  PIN rD[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 0.000 430.640 4.000 ;
    END
  END rD[7]
  PIN rD[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 0.000 438.480 4.000 ;
    END
  END rD[8]
  PIN rD[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 0.000 446.320 4.000 ;
    END
  END rD[9]
  PIN rS[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 0.000 109.200 4.000 ;
    END
  END rS[0]
  PIN rS[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 4.000 ;
    END
  END rS[10]
  PIN rS[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END rS[11]
  PIN rS[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 0.000 203.280 4.000 ;
    END
  END rS[12]
  PIN rS[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 0.000 211.120 4.000 ;
    END
  END rS[13]
  PIN rS[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END rS[14]
  PIN rS[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END rS[15]
  PIN rS[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 0.000 234.640 4.000 ;
    END
  END rS[16]
  PIN rS[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 0.000 242.480 4.000 ;
    END
  END rS[17]
  PIN rS[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 4.000 ;
    END
  END rS[18]
  PIN rS[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 0.000 258.160 4.000 ;
    END
  END rS[19]
  PIN rS[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 4.000 ;
    END
  END rS[1]
  PIN rS[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 0.000 266.000 4.000 ;
    END
  END rS[20]
  PIN rS[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 0.000 273.840 4.000 ;
    END
  END rS[21]
  PIN rS[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 0.000 281.680 4.000 ;
    END
  END rS[22]
  PIN rS[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 0.000 289.520 4.000 ;
    END
  END rS[23]
  PIN rS[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 0.000 297.360 4.000 ;
    END
  END rS[24]
  PIN rS[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.640 0.000 305.200 4.000 ;
    END
  END rS[25]
  PIN rS[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 0.000 313.040 4.000 ;
    END
  END rS[26]
  PIN rS[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 0.000 320.880 4.000 ;
    END
  END rS[27]
  PIN rS[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 0.000 328.720 4.000 ;
    END
  END rS[28]
  PIN rS[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 0.000 336.560 4.000 ;
    END
  END rS[29]
  PIN rS[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END rS[2]
  PIN rS[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 0.000 344.400 4.000 ;
    END
  END rS[30]
  PIN rS[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 0.000 352.240 4.000 ;
    END
  END rS[31]
  PIN rS[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 0.000 132.720 4.000 ;
    END
  END rS[3]
  PIN rS[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 4.000 ;
    END
  END rS[4]
  PIN rS[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 0.000 148.400 4.000 ;
    END
  END rS[5]
  PIN rS[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 4.000 ;
    END
  END rS[6]
  PIN rS[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 0.000 164.080 4.000 ;
    END
  END rS[7]
  PIN rS[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END rS[8]
  PIN rS[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 0.000 179.760 4.000 ;
    END
  END rS[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 784.300 ;
    END
  END vss
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 0.000 367.920 4.000 ;
    END
  END we
  OBS
      LAYER Metal1 ;
        RECT 6.720 4.630 893.200 784.300 ;
      LAYER Metal2 ;
        RECT 4.620 4.300 899.780 784.190 ;
        RECT 4.620 2.330 29.940 4.300 ;
        RECT 31.100 2.330 37.780 4.300 ;
        RECT 38.940 2.330 45.620 4.300 ;
        RECT 46.780 2.330 53.460 4.300 ;
        RECT 54.620 2.330 61.300 4.300 ;
        RECT 62.460 2.330 69.140 4.300 ;
        RECT 70.300 2.330 76.980 4.300 ;
        RECT 78.140 2.330 84.820 4.300 ;
        RECT 85.980 2.330 92.660 4.300 ;
        RECT 93.820 2.330 100.500 4.300 ;
        RECT 101.660 2.330 108.340 4.300 ;
        RECT 109.500 2.330 116.180 4.300 ;
        RECT 117.340 2.330 124.020 4.300 ;
        RECT 125.180 2.330 131.860 4.300 ;
        RECT 133.020 2.330 139.700 4.300 ;
        RECT 140.860 2.330 147.540 4.300 ;
        RECT 148.700 2.330 155.380 4.300 ;
        RECT 156.540 2.330 163.220 4.300 ;
        RECT 164.380 2.330 171.060 4.300 ;
        RECT 172.220 2.330 178.900 4.300 ;
        RECT 180.060 2.330 186.740 4.300 ;
        RECT 187.900 2.330 194.580 4.300 ;
        RECT 195.740 2.330 202.420 4.300 ;
        RECT 203.580 2.330 210.260 4.300 ;
        RECT 211.420 2.330 218.100 4.300 ;
        RECT 219.260 2.330 225.940 4.300 ;
        RECT 227.100 2.330 233.780 4.300 ;
        RECT 234.940 2.330 241.620 4.300 ;
        RECT 242.780 2.330 249.460 4.300 ;
        RECT 250.620 2.330 257.300 4.300 ;
        RECT 258.460 2.330 265.140 4.300 ;
        RECT 266.300 2.330 272.980 4.300 ;
        RECT 274.140 2.330 280.820 4.300 ;
        RECT 281.980 2.330 288.660 4.300 ;
        RECT 289.820 2.330 296.500 4.300 ;
        RECT 297.660 2.330 304.340 4.300 ;
        RECT 305.500 2.330 312.180 4.300 ;
        RECT 313.340 2.330 320.020 4.300 ;
        RECT 321.180 2.330 327.860 4.300 ;
        RECT 329.020 2.330 335.700 4.300 ;
        RECT 336.860 2.330 343.540 4.300 ;
        RECT 344.700 2.330 351.380 4.300 ;
        RECT 352.540 2.330 359.220 4.300 ;
        RECT 360.380 2.330 367.060 4.300 ;
        RECT 368.220 2.330 374.900 4.300 ;
        RECT 376.060 2.330 382.740 4.300 ;
        RECT 383.900 2.330 390.580 4.300 ;
        RECT 391.740 2.330 398.420 4.300 ;
        RECT 399.580 2.330 406.260 4.300 ;
        RECT 407.420 2.330 414.100 4.300 ;
        RECT 415.260 2.330 421.940 4.300 ;
        RECT 423.100 2.330 429.780 4.300 ;
        RECT 430.940 2.330 437.620 4.300 ;
        RECT 438.780 2.330 445.460 4.300 ;
        RECT 446.620 2.330 453.300 4.300 ;
        RECT 454.460 2.330 461.140 4.300 ;
        RECT 462.300 2.330 468.980 4.300 ;
        RECT 470.140 2.330 476.820 4.300 ;
        RECT 477.980 2.330 484.660 4.300 ;
        RECT 485.820 2.330 492.500 4.300 ;
        RECT 493.660 2.330 500.340 4.300 ;
        RECT 501.500 2.330 508.180 4.300 ;
        RECT 509.340 2.330 516.020 4.300 ;
        RECT 517.180 2.330 523.860 4.300 ;
        RECT 525.020 2.330 531.700 4.300 ;
        RECT 532.860 2.330 539.540 4.300 ;
        RECT 540.700 2.330 547.380 4.300 ;
        RECT 548.540 2.330 555.220 4.300 ;
        RECT 556.380 2.330 563.060 4.300 ;
        RECT 564.220 2.330 570.900 4.300 ;
        RECT 572.060 2.330 578.740 4.300 ;
        RECT 579.900 2.330 586.580 4.300 ;
        RECT 587.740 2.330 594.420 4.300 ;
        RECT 595.580 2.330 602.260 4.300 ;
        RECT 603.420 2.330 610.100 4.300 ;
        RECT 611.260 2.330 617.940 4.300 ;
        RECT 619.100 2.330 625.780 4.300 ;
        RECT 626.940 2.330 633.620 4.300 ;
        RECT 634.780 2.330 641.460 4.300 ;
        RECT 642.620 2.330 649.300 4.300 ;
        RECT 650.460 2.330 657.140 4.300 ;
        RECT 658.300 2.330 664.980 4.300 ;
        RECT 666.140 2.330 672.820 4.300 ;
        RECT 673.980 2.330 680.660 4.300 ;
        RECT 681.820 2.330 688.500 4.300 ;
        RECT 689.660 2.330 696.340 4.300 ;
        RECT 697.500 2.330 704.180 4.300 ;
        RECT 705.340 2.330 712.020 4.300 ;
        RECT 713.180 2.330 719.860 4.300 ;
        RECT 721.020 2.330 727.700 4.300 ;
        RECT 728.860 2.330 735.540 4.300 ;
        RECT 736.700 2.330 743.380 4.300 ;
        RECT 744.540 2.330 751.220 4.300 ;
        RECT 752.380 2.330 759.060 4.300 ;
        RECT 760.220 2.330 766.900 4.300 ;
        RECT 768.060 2.330 774.740 4.300 ;
        RECT 775.900 2.330 782.580 4.300 ;
        RECT 783.740 2.330 790.420 4.300 ;
        RECT 791.580 2.330 798.260 4.300 ;
        RECT 799.420 2.330 806.100 4.300 ;
        RECT 807.260 2.330 813.940 4.300 ;
        RECT 815.100 2.330 821.780 4.300 ;
        RECT 822.940 2.330 829.620 4.300 ;
        RECT 830.780 2.330 837.460 4.300 ;
        RECT 838.620 2.330 845.300 4.300 ;
        RECT 846.460 2.330 853.140 4.300 ;
        RECT 854.300 2.330 860.980 4.300 ;
        RECT 862.140 2.330 868.820 4.300 ;
        RECT 869.980 2.330 899.780 4.300 ;
      LAYER Metal3 ;
        RECT 4.570 2.380 899.830 784.140 ;
      LAYER Metal4 ;
        RECT 10.780 19.130 21.940 715.590 ;
        RECT 24.140 19.130 98.740 715.590 ;
        RECT 100.940 19.130 175.540 715.590 ;
        RECT 177.740 19.130 252.340 715.590 ;
        RECT 254.540 19.130 329.140 715.590 ;
        RECT 331.340 19.130 405.940 715.590 ;
        RECT 408.140 19.130 482.740 715.590 ;
        RECT 484.940 19.130 559.540 715.590 ;
        RECT 561.740 19.130 636.340 715.590 ;
        RECT 638.540 19.130 713.140 715.590 ;
        RECT 715.340 19.130 789.940 715.590 ;
        RECT 792.140 19.130 866.740 715.590 ;
        RECT 868.940 19.130 881.300 715.590 ;
  END
END minimax_rf
END LIBRARY

